/*  This file is part of JTCORES.
    JTCORES program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTCORES program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTCORES.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 23-8-2025 */

module jtrungun_dim(
    input             rst,   clk, pxl_cen,
                      lhbl, lvbl,

    output     [11:1] pal_addr,
    input      [15:0] pal_dout,

    input      [15:0] pxl,

    output     [ 7:0] red,
    output     [ 7:0] green,
    output     [ 7:0] blue
);

reg  [23:0] bgr;
wire [ 7:0] r8, b8, g8;
wire        shad;

assign {blue,green,red} = (lvbl & lhbl ) ? bgr : 24'd0;
assign pal_addr = pxl[11:1];

function [7:0] conv58(input [4:0] cin );
begin
    conv58 = {cin, cin[4-:3]};
end
endfunction

assign { b8, g8, r8 } = {conv58(pal_dout[10+:5]),conv58(pal_dout[5+:5]),conv58(pal_dout[0+:5])};
assign shad = pxl[0];

always @(posedge clk) begin
    if( rst ) begin
        bgr   <= 0;
    end else begin
        if( pxl_cen ) bgr <= ~shad ? { b8, g8, r8 } : { b8>>1, g8>>1, r8>>1 };
    end
end

endmodule