../../1942/hdl/1942.vh