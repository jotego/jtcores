/* verilator lint_off UNOPTFLAT */

module vlm5030_delay_21
  (input  i_clk_base,
   input  i_clk_val,
   input  i_clk_rise,
   input  i_clk_fall,
   input  i_in,
   output o_out);
  wire [3:0] n20773_o;
  reg [30:0] delay_p_cnt;
  reg delay_p_inq;
  wire n20783_o;
  wire n20785_o;
  wire n20787_o;
  wire [31:0] n20788_o;
  wire n20790_o;
  wire [31:0] n20791_o;
  wire [31:0] n20793_o;
  wire [30:0] n20794_o;
  wire n20795_o;
  wire [30:0] n20796_o;
  wire n20797_o;
  wire [30:0] n20799_o;
  wire [30:0] n20805_o;
  reg [30:0] n20806_q;
  wire n20807_o;
  wire n20808_o;
  reg n20809_q;
  wire n20810_o;
  reg n20811_q;
  assign o_out = n20811_q;
  /* clock_functions_pack.vhd:57:15  */
  assign n20773_o = {i_clk_fall, i_clk_rise, i_clk_val, i_clk_base};
  /* vlm5030_subcircuits.vhd:129:14  */
  always @*
    delay_p_cnt = n20806_q; // (isignal)
  initial
    delay_p_cnt = 31'b0000000000000000000000000000000;
  /* vlm5030_subcircuits.vhd:130:14  */
  always @*
    delay_p_inq = n20809_q; // (isignal)
  initial
    delay_p_inq = 1'b0;
  /* clock_functions_pack.vhd:36:12  */
  assign n20783_o = n20773_o[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n20785_o = n20773_o[2];
  /* vlm5030_subcircuits.vhd:133:15  */
  assign n20787_o = i_in != delay_p_inq;
  /* vlm5030_subcircuits.vhd:137:16  */
  assign n20788_o = {1'b0, delay_p_cnt};  //  uext
  /* vlm5030_subcircuits.vhd:137:16  */
  assign n20790_o = $signed(n20788_o) > $signed(32'b00000000000000000000000000000000);
  /* vlm5030_subcircuits.vhd:138:22  */
  assign n20791_o = {1'b0, delay_p_cnt};  //  uext
  /* vlm5030_subcircuits.vhd:138:22  */
  assign n20793_o = n20791_o - 32'b00000000000000000000000000000001;
  /* vlm5030_subcircuits.vhd:138:11  */
  assign n20794_o = n20793_o[30:0];  // trunc
  /* vlm5030_subcircuits.vhd:137:9  */
  assign n20795_o = n20790_o ? n20811_q : i_in;
  /* vlm5030_subcircuits.vhd:137:9  */
  assign n20796_o = n20790_o ? n20794_o : delay_p_cnt;
  /* vlm5030_subcircuits.vhd:133:7  */
  assign n20797_o = n20787_o ? n20811_q : n20795_o;
  /* vlm5030_subcircuits.vhd:133:7  */
  assign n20799_o = n20787_o ? 31'b0000000000000000000000000010011 : n20796_o;
  /* vlm5030_subcircuits.vhd:132:5  */
  assign n20805_o = n20785_o ? n20799_o : delay_p_cnt;
  /* vlm5030_subcircuits.vhd:132:5  */
  always @(posedge n20783_o)
    n20806_q <= n20805_o;
  initial
    n20806_q = 31'b0000000000000000000000000000000;
  /* vlm5030_subcircuits.vhd:132:5  */
  assign n20807_o = n20785_o & n20787_o;
  /* vlm5030_subcircuits.vhd:132:5  */
  assign n20808_o = n20807_o ? i_in : delay_p_inq;
  /* vlm5030_subcircuits.vhd:132:5  */
  always @(posedge n20783_o)
    n20809_q <= n20808_o;
  initial
    n20809_q = 1'b0;
  /* vlm5030_subcircuits.vhd:132:5  */
  assign n20810_o = n20785_o ? n20797_o : n20811_q;
  /* vlm5030_subcircuits.vhd:132:5  */
  always @(posedge n20783_o)
    n20811_q <= n20810_o;
endmodule

module vlm5030_srlatch
  (input  i_clk,
   input  i_res,
   input  i_set,
   output o_q);
  reg q;
  wire n20767_o;
  wire n20769_o;
  reg n20772_q;
  assign o_q = q;
  /* vlm5030_subcircuits.vhd:37:10  */
  always @*
    q = n20772_q; // (isignal)
  initial
    q = 1'b0;
  /* vlm5030_subcircuits.vhd:45:7  */
  assign n20767_o = i_set ? 1'b1 : q;
  /* vlm5030_subcircuits.vhd:43:7  */
  assign n20769_o = i_res ? 1'b0 : n20767_o;
  /* vlm5030_subcircuits.vhd:42:5  */
  always @(posedge i_clk)
    n20772_q <= n20769_o;
  initial
    n20772_q = 1'b0;
endmodule

module vlm5030_delay_4
  (input  i_clk_base,
   input  i_clk_val,
   input  i_clk_rise,
   input  i_clk_fall,
   input  i_in,
   output o_out);
  wire [3:0] n20722_o;
  reg [30:0] delay_p_cnt;
  reg delay_p_inq;
  wire n20732_o;
  wire n20734_o;
  wire n20736_o;
  wire [31:0] n20737_o;
  wire n20739_o;
  wire [31:0] n20740_o;
  wire [31:0] n20742_o;
  wire [30:0] n20743_o;
  wire n20744_o;
  wire [30:0] n20745_o;
  wire n20746_o;
  wire [30:0] n20748_o;
  wire [30:0] n20754_o;
  reg [30:0] n20755_q;
  wire n20756_o;
  wire n20757_o;
  reg n20758_q;
  wire n20759_o;
  reg n20760_q;
  assign o_out = n20760_q;
  /* clock_functions_pack.vhd:51:14  */
  assign n20722_o = {i_clk_fall, i_clk_rise, i_clk_val, i_clk_base};
  /* vlm5030_subcircuits.vhd:129:14  */
  always @*
    delay_p_cnt = n20755_q; // (isignal)
  initial
    delay_p_cnt = 31'b0000000000000000000000000000000;
  /* vlm5030_subcircuits.vhd:130:14  */
  always @*
    delay_p_inq = n20758_q; // (isignal)
  initial
    delay_p_inq = 1'b0;
  /* vlm5030_gl.vhd:1779:14  */
  assign n20732_o = n20722_o[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n20734_o = n20722_o[2];
  /* vlm5030_subcircuits.vhd:133:15  */
  assign n20736_o = i_in != delay_p_inq;
  /* vlm5030_subcircuits.vhd:137:16  */
  assign n20737_o = {1'b0, delay_p_cnt};  //  uext
  /* vlm5030_subcircuits.vhd:137:16  */
  assign n20739_o = $signed(n20737_o) > $signed(32'b00000000000000000000000000000000);
  /* vlm5030_subcircuits.vhd:138:22  */
  assign n20740_o = {1'b0, delay_p_cnt};  //  uext
  /* vlm5030_subcircuits.vhd:138:22  */
  assign n20742_o = n20740_o - 32'b00000000000000000000000000000001;
  /* vlm5030_subcircuits.vhd:138:11  */
  assign n20743_o = n20742_o[30:0];  // trunc
  /* vlm5030_subcircuits.vhd:137:9  */
  assign n20744_o = n20739_o ? n20760_q : i_in;
  /* vlm5030_subcircuits.vhd:137:9  */
  assign n20745_o = n20739_o ? n20743_o : delay_p_cnt;
  /* vlm5030_subcircuits.vhd:133:7  */
  assign n20746_o = n20736_o ? n20760_q : n20744_o;
  /* vlm5030_subcircuits.vhd:133:7  */
  assign n20748_o = n20736_o ? 31'b0000000000000000000000000000010 : n20745_o;
  /* vlm5030_subcircuits.vhd:132:5  */
  assign n20754_o = n20734_o ? n20748_o : delay_p_cnt;
  /* vlm5030_subcircuits.vhd:132:5  */
  always @(posedge n20732_o)
    n20755_q <= n20754_o;
  initial
    n20755_q = 31'b0000000000000000000000000000000;
  /* vlm5030_subcircuits.vhd:132:5  */
  assign n20756_o = n20734_o & n20736_o;
  /* vlm5030_subcircuits.vhd:132:5  */
  assign n20757_o = n20756_o ? i_in : delay_p_inq;
  /* vlm5030_subcircuits.vhd:132:5  */
  always @(posedge n20732_o)
    n20758_q <= n20757_o;
  initial
    n20758_q = 1'b0;
  /* vlm5030_subcircuits.vhd:132:5  */
  assign n20759_o = n20734_o ? n20746_o : n20760_q;
  /* vlm5030_subcircuits.vhd:132:5  */
  always @(posedge n20732_o)
    n20760_q <= n20759_o;
endmodule

module vlm5030_delay_inv_4
  (input  i_clk_base,
   input  i_clk_val,
   input  i_clk_rise,
   input  i_clk_fall,
   input  i_in,
   output o_out);
  wire [3:0] n20678_o;
  wire outq;
  reg [30:0] delay_p_cnt;
  reg delay_p_inq;
  wire n20688_o;
  wire n20690_o;
  wire n20692_o;
  wire n20694_o;
  wire [31:0] n20695_o;
  wire n20697_o;
  wire [31:0] n20698_o;
  wire [31:0] n20700_o;
  wire [30:0] n20701_o;
  wire n20702_o;
  wire [30:0] n20703_o;
  wire n20704_o;
  wire [30:0] n20706_o;
  wire [30:0] n20712_o;
  reg [30:0] n20713_q;
  wire n20714_o;
  wire n20715_o;
  reg n20716_q;
  wire n20718_o;
  wire n20719_o;
  wire n20720_o;
  reg n20721_q;
  assign o_out = n20718_o;
  assign n20678_o = {i_clk_fall, i_clk_rise, i_clk_val, i_clk_base};
  /* vlm5030_subcircuits.vhd:177:10  */
  assign outq = n20721_q; // (signal)
  /* vlm5030_subcircuits.vhd:181:14  */
  always @*
    delay_p_cnt = n20713_q; // (isignal)
  initial
    delay_p_cnt = 31'b0000000000000000000000000000000;
  /* vlm5030_subcircuits.vhd:182:14  */
  always @*
    delay_p_inq = n20716_q; // (isignal)
  initial
    delay_p_inq = 1'b0;
  /* clock_functions_pack.vhd:36:12  */
  assign n20688_o = n20678_o[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n20690_o = n20678_o[2];
  /* vlm5030_subcircuits.vhd:185:15  */
  assign n20692_o = i_in != delay_p_inq;
  /* vlm5030_subcircuits.vhd:188:9  */
  assign n20694_o = i_in ? 1'b1 : outq;
  /* vlm5030_subcircuits.vhd:192:16  */
  assign n20695_o = {1'b0, delay_p_cnt};  //  uext
  /* vlm5030_subcircuits.vhd:192:16  */
  assign n20697_o = $signed(n20695_o) > $signed(32'b00000000000000000000000000000000);
  /* vlm5030_subcircuits.vhd:193:22  */
  assign n20698_o = {1'b0, delay_p_cnt};  //  uext
  /* vlm5030_subcircuits.vhd:193:22  */
  assign n20700_o = n20698_o - 32'b00000000000000000000000000000001;
  /* vlm5030_subcircuits.vhd:193:11  */
  assign n20701_o = n20700_o[30:0];  // trunc
  /* vlm5030_subcircuits.vhd:192:9  */
  assign n20702_o = n20697_o ? outq : i_in;
  /* vlm5030_subcircuits.vhd:192:9  */
  assign n20703_o = n20697_o ? n20701_o : delay_p_cnt;
  /* vlm5030_subcircuits.vhd:185:7  */
  assign n20704_o = n20692_o ? n20694_o : n20702_o;
  /* vlm5030_subcircuits.vhd:185:7  */
  assign n20706_o = n20692_o ? 31'b0000000000000000000000000000010 : n20703_o;
  /* vlm5030_subcircuits.vhd:184:5  */
  assign n20712_o = n20690_o ? n20706_o : delay_p_cnt;
  /* vlm5030_subcircuits.vhd:184:5  */
  always @(posedge n20688_o)
    n20713_q <= n20712_o;
  initial
    n20713_q = 31'b0000000000000000000000000000000;
  /* vlm5030_subcircuits.vhd:184:5  */
  assign n20714_o = n20690_o & n20692_o;
  /* vlm5030_subcircuits.vhd:184:5  */
  assign n20715_o = n20714_o ? i_in : delay_p_inq;
  /* vlm5030_subcircuits.vhd:184:5  */
  always @(posedge n20688_o)
    n20716_q <= n20715_o;
  initial
    n20716_q = 1'b0;
  /* vlm5030_subcircuits.vhd:201:16  */
  assign n20718_o = i_in ? 1'b0 : n20719_o;
  /* vlm5030_subcircuits.vhd:201:37  */
  assign n20719_o = ~outq;
  /* vlm5030_subcircuits.vhd:184:5  */
  assign n20720_o = n20690_o ? n20704_o : outq;
  /* vlm5030_subcircuits.vhd:184:5  */
  always @(posedge n20688_o)
    n20721_q <= n20720_o;
endmodule

module vlm5030_delay_inv_2
  (input  i_clk_base,
   input  i_clk_val,
   input  i_clk_rise,
   input  i_clk_fall,
   input  i_in,
   output o_out);
  wire [3:0] n20634_o;
  wire outq;
  reg [30:0] delay_p_cnt;
  reg delay_p_inq;
  wire n20644_o;
  wire n20646_o;
  wire n20648_o;
  wire n20650_o;
  wire [31:0] n20651_o;
  wire n20653_o;
  wire [31:0] n20654_o;
  wire [31:0] n20656_o;
  wire [30:0] n20657_o;
  wire n20658_o;
  wire [30:0] n20659_o;
  wire n20660_o;
  wire [30:0] n20662_o;
  wire [30:0] n20668_o;
  reg [30:0] n20669_q;
  wire n20670_o;
  wire n20671_o;
  reg n20672_q;
  wire n20674_o;
  wire n20675_o;
  wire n20676_o;
  reg n20677_q;
  assign o_out = n20674_o;
  assign n20634_o = {i_clk_fall, i_clk_rise, i_clk_val, i_clk_base};
  /* vlm5030_subcircuits.vhd:177:10  */
  assign outq = n20677_q; // (signal)
  /* vlm5030_subcircuits.vhd:181:14  */
  always @*
    delay_p_cnt = n20669_q; // (isignal)
  initial
    delay_p_cnt = 31'b0000000000000000000000000000000;
  /* vlm5030_subcircuits.vhd:182:14  */
  always @*
    delay_p_inq = n20672_q; // (isignal)
  initial
    delay_p_inq = 1'b0;
  assign n20644_o = n20634_o[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n20646_o = n20634_o[2];
  /* vlm5030_subcircuits.vhd:185:15  */
  assign n20648_o = i_in != delay_p_inq;
  /* vlm5030_subcircuits.vhd:188:9  */
  assign n20650_o = i_in ? 1'b1 : outq;
  /* vlm5030_subcircuits.vhd:192:16  */
  assign n20651_o = {1'b0, delay_p_cnt};  //  uext
  /* vlm5030_subcircuits.vhd:192:16  */
  assign n20653_o = $signed(n20651_o) > $signed(32'b00000000000000000000000000000000);
  /* vlm5030_subcircuits.vhd:193:22  */
  assign n20654_o = {1'b0, delay_p_cnt};  //  uext
  /* vlm5030_subcircuits.vhd:193:22  */
  assign n20656_o = n20654_o - 32'b00000000000000000000000000000001;
  /* vlm5030_subcircuits.vhd:193:11  */
  assign n20657_o = n20656_o[30:0];  // trunc
  /* vlm5030_subcircuits.vhd:192:9  */
  assign n20658_o = n20653_o ? outq : i_in;
  /* vlm5030_subcircuits.vhd:192:9  */
  assign n20659_o = n20653_o ? n20657_o : delay_p_cnt;
  /* vlm5030_subcircuits.vhd:185:7  */
  assign n20660_o = n20648_o ? n20650_o : n20658_o;
  /* vlm5030_subcircuits.vhd:185:7  */
  assign n20662_o = n20648_o ? 31'b0000000000000000000000000000000 : n20659_o;
  /* vlm5030_subcircuits.vhd:184:5  */
  assign n20668_o = n20646_o ? n20662_o : delay_p_cnt;
  /* vlm5030_subcircuits.vhd:184:5  */
  always @(posedge n20644_o)
    n20669_q <= n20668_o;
  initial
    n20669_q = 31'b0000000000000000000000000000000;
  /* vlm5030_subcircuits.vhd:184:5  */
  assign n20670_o = n20646_o & n20648_o;
  /* vlm5030_subcircuits.vhd:184:5  */
  assign n20671_o = n20670_o ? i_in : delay_p_inq;
  /* vlm5030_subcircuits.vhd:184:5  */
  always @(posedge n20644_o)
    n20672_q <= n20671_o;
  initial
    n20672_q = 1'b0;
  /* vlm5030_subcircuits.vhd:201:16  */
  assign n20674_o = i_in ? 1'b0 : n20675_o;
  /* vlm5030_subcircuits.vhd:201:37  */
  assign n20675_o = ~outq;
  /* vlm5030_subcircuits.vhd:184:5  */
  assign n20676_o = n20646_o ? n20660_o : outq;
  /* vlm5030_subcircuits.vhd:184:5  */
  always @(posedge n20644_o)
    n20677_q <= n20676_o;
endmodule

module vlm5030_srlatchclk
  (input  i_clk_base,
   input  i_clk_val,
   input  i_clk_rise,
   input  i_clk_fall,
   input  i_res_base,
   input  i_res_val,
   input  i_res_rise,
   input  i_res_fall,
   input  i_set_base,
   input  i_set_val,
   input  i_set_rise,
   input  i_set_fall,
   output o_q_base,
   output o_q_val,
   output o_q_rise,
   output o_q_fall);
  wire [3:0] n20597_o;
  wire [3:0] n20598_o;
  wire [3:0] n20599_o;
  wire n20601_o;
  wire n20602_o;
  wire n20603_o;
  wire n20604_o;
  reg q;
  wire n20613_o;
  wire n20615_o;
  wire n20617_o;
  wire n20618_o;
  wire n20620_o;
  wire n20622_o;
  wire n20625_o;
  wire n20626_o;
  wire n20627_o;
  wire n20628_o;
  wire n20629_o;
  wire n20630_o;
  wire [3:0] n20631_o;
  wire n20632_o;
  reg n20633_q;
  assign o_q_base = n20601_o;
  assign o_q_val = n20602_o;
  assign o_q_rise = n20603_o;
  assign o_q_fall = n20604_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20597_o = {i_clk_fall, i_clk_rise, i_clk_val, i_clk_base};
  /* vlm5030_pack.vhd:27:13  */
  assign n20598_o = {i_res_fall, i_res_rise, i_res_val, i_res_base};
  /* vlm5030_pack.vhd:27:13  */
  assign n20599_o = {i_set_fall, i_set_rise, i_set_val, i_set_base};
  /* vlm5030_pack.vhd:27:13  */
  assign n20601_o = n20631_o[0];
  assign n20602_o = n20631_o[1];
  /* vlm5030_pack.vhd:46:14  */
  assign n20603_o = n20631_o[2];
  assign n20604_o = n20631_o[3];
  /* vlm5030_subcircuits.vhd:77:10  */
  always @*
    q = n20633_q; // (isignal)
  initial
    q = 1'b0;
  /* vlm5030_pack.vhd:27:13  */
  assign n20613_o = n20597_o[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n20615_o = n20597_o[2];
  /* vlm5030_subcircuits.vhd:83:16  */
  assign n20617_o = n20598_o[1];
  /* vlm5030_subcircuits.vhd:85:19  */
  assign n20618_o = n20599_o[1];
  /* vlm5030_subcircuits.vhd:85:7  */
  assign n20620_o = n20618_o ? 1'b1 : q;
  /* vlm5030_subcircuits.vhd:83:7  */
  assign n20622_o = n20617_o ? 1'b0 : n20620_o;
  /* vlm5030_subcircuits.vhd:91:25  */
  assign n20625_o = n20597_o[0];
  /* vlm5030_subcircuits.vhd:93:19  */
  assign n20626_o = ~q;
  /* vlm5030_subcircuits.vhd:93:35  */
  assign n20627_o = n20599_o[1];
  /* vlm5030_subcircuits.vhd:93:25  */
  assign n20628_o = n20626_o & n20627_o;
  /* vlm5030_subcircuits.vhd:94:35  */
  assign n20629_o = n20598_o[1];
  /* vlm5030_subcircuits.vhd:94:25  */
  assign n20630_o = q & n20629_o;
  assign n20631_o = {n20630_o, n20628_o, q, n20625_o};
  /* vlm5030_subcircuits.vhd:82:5  */
  assign n20632_o = n20615_o ? n20622_o : q;
  /* vlm5030_subcircuits.vhd:82:5  */
  always @(posedge n20613_o)
    n20633_q <= n20632_o;
  initial
    n20633_q = 1'b0;
endmodule

module vlm5030_gl
  (input  i_clk,
   input  i_oscen,
   input  i_rst,
   input  i_start,
   input  i_vcu,
   input  i_vref,
   input  i_tst1,
   input  i_tst3,
   input  [7:0] i_d,
   output o_tst2,
   output o_tst4,
   output [15:0] o_a,
   output o_me_l,
   output o_mte,
   output o_bsy,
   output [5:0] o_dao,
   output [9:0] o_audio);
  wire [3:0] osc;
  localparam [3:0] n8_o = 4'b0000;
  reg [3:0] clk2;
  wire [3:0] nclk2;
  wire rst;
  wire [7:0] dq;
  wire maskdq53;
  wire starttst;
  wire tststopclk2;
  wire tstend2id;
  wire tstend2ie;
  wire tstenid2a;
  wire tstenie2a;
  wire tstenctrl2a;
  wire tstenie2dac;
  reg [10:0] clk2divq;
  wire [3:0] c2d0;
  wire [3:0] c2d1;
  wire [3:0] c2d3;
  wire [3:0] c2d4;
  wire [3:0] c2d5;
  wire [3:0] c2d6;
  wire [3:0] c2d7;
  wire [3:0] c2d8;
  wire [3:0] c2d9;
  wire [3:0] c2d10;
  wire [3:0] c2d5fin;
  wire [3:0] c2d7fin;
  wire [3:0] nc2d7fin;
  wire [3:0] c2d9fin;
  wire [3:0] nc2d9fin;
  wire [3:0] clk2gd5;
  wire [3:0] nc2d1;
  wire [3:0] nc2d6;
  wire [3:0] nc2d8;
  wire [3:0] nc2d10;
  wire [3:0] c2d3gated;
  wire fsromevalout;
  wire [13:0] fsromdo;
  wire fsromnorhigh;
  wire fsromnorlow;
  wire [3:0] clk2ctrl;
  wire ncen1;
  wire cen3;
  wire eaoen;
  reg xromdo7nq;
  wire xromdo7q;
  wire [36:0] xromdo;
  wire [4:0] yromdo;
  wire c2d3gate;
  wire cntdn0;
  reg [7:0] dinalq;
  wire [15:0] aq;
  wire startrise;
  wire [3:0] clkcntdn;
  wire ncntdnload;
  wire ncntdn;
  wire eavcu;
  wire ealatchh;
  wire neaload;
  wire eainc;
  wire clrdinal;
  wire clkdin;
  wire nvcufinal;
  wire vcufinal12;
  wire nbsy;
  wire me;
  wire rflatchwen;
  wire asshift2;
  wire updtpitch;
  wire enrf2id;
  wire [3:0] clkksa;
  wire ensum2id;
  wire [3:0] clk2ena;
  wire [3:0] clk2enb;
  wire rstdel;
  wire [4:0] ksa;
  wire [9:0] nkdo;
  wire [9:0] rfdo;
  wire rfdo97zero;
  wire [9:0] nid;
  wire [9:0] assum;
  wire [11:0] nie;
  wire [7:0] idlat;
  wire idlatall1;
  wire enidlinv2id;
  wire enidl2ie;
  wire enidlinv2ie;
  wire pitchoverflow;
  wire [3:0] enpitchlat;
  wire enmem02id;
  wire [9:0] nmem0do;
  wire [9:0] mem0do;
  wire enmem12ie;
  wire [11:0] mem1do2ie;
  wire enmem22ie;
  wire [11:0] mem2do2ie;
  wire [11:0] ieregdrv;
  wire [11:0] ieregdrv4ie;
  wire [3:0] ieregload;
  wire enieregfa2ie;
  wire [3:0] c2d10xr9;
  wire enie2a;
  wire [11:0] ieaddrreg;
  wire pitchmod;
  wire random;
  wire pwmsr;
  wire [3:0] n14_o;
  wire n17_o;
  wire n22_o;
  wire n23_o;
  wire n24_o;
  wire n25_o;
  wire n26_o;
  wire n27_o;
  wire n28_o;
  wire n29_o;
  wire n30_o;
  wire [3:0] n31_o;
  wire n36_o;
  wire n37_o;
  wire n38_o;
  wire n39_o;
  wire n40_o;
  wire n41_o;
  wire n42_o;
  wire n43_o;
  wire n44_o;
  wire [3:0] n45_o;
  wire n49_o;
  wire n54_o;
  wire n55_o;
  wire n56_o;
  wire n57_o;
  wire n58_o;
  wire n59_o;
  wire n60_o;
  wire n61_o;
  wire n62_o;
  wire [3:0] n63_o;
  wire n68_o;
  wire n69_o;
  wire n70_o;
  wire n71_o;
  wire n72_o;
  wire n73_o;
  wire n74_o;
  wire n75_o;
  wire n76_o;
  wire [3:0] n77_o;
  wire n78_o;
  wire n79_o;
  wire n84_o;
  wire n85_o;
  wire n86_o;
  wire n87_o;
  wire n88_o;
  wire n89_o;
  wire n90_o;
  wire n91_o;
  wire n92_o;
  wire [3:0] n93_o;
  reg [7:0] rstdel_block_porcnt;
  reg rstdel_block_npor;
  reg [1:0] rstdel_block_del;
  wire n103_o;
  wire n105_o;
  wire n106_o;
  wire n108_o;
  wire [7:0] n110_o;
  wire n113_o;
  wire n119_o;
  wire n121_o;
  wire n122_o;
  wire n123_o;
  wire n130_o;
  wire n132_o;
  wire n134_o;
  wire [1:0] n135_o;
  wire n138_o;
  wire n139_o;
  wire [7:0] n140_o;
  reg [7:0] n141_q;
  wire n142_o;
  reg n143_q;
  wire [1:0] n144_o;
  reg [1:0] n145_q;
  reg dq_block_rstq;
  wire [3:0] dq_block_rstclk;
  wire [7:0] dq_block_ldq;
  reg dq_block_maskdq53m;
  reg dq_block_maskdq53s;
  wire n150_o;
  wire n154_o;
  wire n155_o;
  wire n156_o;
  wire n157_o;
  wire n158_o;
  wire [3:0] n159_o;
  wire n166_o;
  wire n168_o;
  wire n178_o;
  wire n180_o;
  wire n192_o;
  wire n194_o;
  wire [2:0] n202_o;
  wire [2:0] n203_o;
  wire [1:0] n204_o;
  wire [2:0] n205_o;
  reg n207_q;
  wire [7:0] n208_o;
  reg [7:0] n209_q;
  wire n210_o;
  reg n211_q;
  wire n212_o;
  reg n213_q;
  wire tst_block_ntst1;
  wire tst_block_nstart;
  wire tst_block_nvcu;
  wire tst_block_ntst1vref;
  wire n214_o;
  wire n215_o;
  wire n216_o;
  wire n217_o;
  wire n218_o;
  wire n219_o;
  wire n220_o;
  wire n221_o;
  wire n222_o;
  wire n223_o;
  wire n224_o;
  wire n225_o;
  wire n226_o;
  wire n227_o;
  wire n228_o;
  wire n229_o;
  wire n230_o;
  wire n231_o;
  wire n232_o;
  wire n233_o;
  wire n234_o;
  wire n235_o;
  wire n236_o;
  wire n237_o;
  wire n238_o;
  wire n239_o;
  wire n240_o;
  wire n241_o;
  wire n242_o;
  wire n243_o;
  wire n251_o;
  wire n253_o;
  wire n256_o;
  wire n257_o;
  wire n258_o;
  wire n263_o;
  wire n264_o;
  wire n270_o;
  wire n271_o;
  wire n272_o;
  wire n275_o;
  wire n276_o;
  wire n282_o;
  wire n283_o;
  wire n290_o;
  wire n291_o;
  wire n292_o;
  wire n293_o;
  wire n294_o;
  wire [3:0] n295_o;
  wire clk2div_block_c2qnor;
  wire clk2div_block_feedback;
  wire n303_o;
  wire n305_o;
  wire [9:0] n307_o;
  wire [10:0] n308_o;
  wire [9:0] n312_o;
  wire n318_o;
  wire n320_o;
  wire n322_o;
  wire n323_o;
  wire n324_o;
  wire n325_o;
  wire n326_o;
  wire n327_o;
  wire n328_o;
  wire n329_o;
  wire n330_o;
  wire n331_o;
  wire n332_o;
  wire n333_o;
  wire n334_o;
  wire n335_o;
  wire n336_o;
  wire n337_o;
  wire n338_o;
  wire n339_o;
  wire n340_o;
  wire n342_o;
  wire n344_o;
  wire n349_o;
  wire n350_o;
  wire n351_o;
  wire n352_o;
  wire n353_o;
  wire n354_o;
  wire n355_o;
  wire n356_o;
  wire n357_o;
  wire [3:0] n358_o;
  wire n360_o;
  wire n361_o;
  wire n366_o;
  wire n367_o;
  wire n368_o;
  wire n369_o;
  wire n370_o;
  wire n371_o;
  wire n372_o;
  wire n373_o;
  wire n374_o;
  wire [3:0] n375_o;
  wire n377_o;
  wire n378_o;
  wire n383_o;
  wire n384_o;
  wire n385_o;
  wire n386_o;
  wire n387_o;
  wire n388_o;
  wire n389_o;
  wire n390_o;
  wire n391_o;
  wire [3:0] n392_o;
  wire n394_o;
  wire n395_o;
  wire n400_o;
  wire n401_o;
  wire n402_o;
  wire n403_o;
  wire n404_o;
  wire n405_o;
  wire n406_o;
  wire n407_o;
  wire n408_o;
  wire [3:0] n409_o;
  wire n411_o;
  wire n412_o;
  wire n417_o;
  wire n418_o;
  wire n419_o;
  wire n420_o;
  wire n421_o;
  wire n422_o;
  wire n423_o;
  wire n424_o;
  wire n425_o;
  wire [3:0] n426_o;
  wire n428_o;
  wire n429_o;
  wire n434_o;
  wire n435_o;
  wire n436_o;
  wire n437_o;
  wire n438_o;
  wire n439_o;
  wire n440_o;
  wire n441_o;
  wire n442_o;
  wire [3:0] n443_o;
  wire n445_o;
  wire n446_o;
  wire n451_o;
  wire n452_o;
  wire n453_o;
  wire n454_o;
  wire n455_o;
  wire n456_o;
  wire n457_o;
  wire n458_o;
  wire n459_o;
  wire [3:0] n460_o;
  wire n462_o;
  wire n463_o;
  wire n468_o;
  wire n469_o;
  wire n470_o;
  wire n471_o;
  wire n472_o;
  wire n473_o;
  wire n474_o;
  wire n475_o;
  wire n476_o;
  wire [3:0] n477_o;
  wire n479_o;
  wire n480_o;
  wire n485_o;
  wire n486_o;
  wire n487_o;
  wire n488_o;
  wire n489_o;
  wire n490_o;
  wire n491_o;
  wire n492_o;
  wire n493_o;
  wire [3:0] n494_o;
  wire n496_o;
  wire n497_o;
  wire n502_o;
  wire n503_o;
  wire n504_o;
  wire n505_o;
  wire n506_o;
  wire n507_o;
  wire n508_o;
  wire n509_o;
  wire n510_o;
  wire [3:0] n511_o;
  wire clk2div_block_c2d5fin_b_o_q_base;
  wire clk2div_block_c2d5fin_b_o_q_val;
  wire clk2div_block_c2d5fin_b_o_q_rise;
  wire clk2div_block_c2d5fin_b_o_q_fall;
  wire n512_o;
  wire n513_o;
  wire n514_o;
  wire n515_o;
  wire n516_o;
  wire n517_o;
  wire n518_o;
  wire n519_o;
  wire n520_o;
  wire n521_o;
  wire n522_o;
  wire n523_o;
  wire [3:0] n524_o;
  wire clk2div_block_c2d7fin_b_o_q_base;
  wire clk2div_block_c2d7fin_b_o_q_val;
  wire clk2div_block_c2d7fin_b_o_q_rise;
  wire clk2div_block_c2d7fin_b_o_q_fall;
  wire n526_o;
  wire n527_o;
  wire n528_o;
  wire n529_o;
  wire n530_o;
  wire n531_o;
  wire n532_o;
  wire n533_o;
  wire n534_o;
  wire n535_o;
  wire n536_o;
  wire n537_o;
  wire [3:0] n538_o;
  wire n545_o;
  wire n546_o;
  wire n547_o;
  wire n548_o;
  wire n549_o;
  wire [3:0] n550_o;
  wire clk2div_block_c2d9fin_b_o_q_base;
  wire clk2div_block_c2d9fin_b_o_q_val;
  wire clk2div_block_c2d9fin_b_o_q_rise;
  wire clk2div_block_c2d9fin_b_o_q_fall;
  wire n551_o;
  wire n552_o;
  wire n553_o;
  wire n554_o;
  wire n555_o;
  wire n556_o;
  wire n557_o;
  wire n558_o;
  wire n559_o;
  wire n560_o;
  wire n561_o;
  wire n562_o;
  wire [3:0] n563_o;
  wire n570_o;
  wire n571_o;
  wire n572_o;
  wire n573_o;
  wire n574_o;
  wire [3:0] n575_o;
  wire n582_o;
  wire n583_o;
  wire n584_o;
  wire n585_o;
  wire n586_o;
  wire n587_o;
  wire n588_o;
  wire n589_o;
  wire n590_o;
  wire n591_o;
  wire n592_o;
  wire n593_o;
  wire n594_o;
  wire n595_o;
  wire n596_o;
  wire n597_o;
  wire n598_o;
  wire n599_o;
  wire n600_o;
  wire n601_o;
  wire n602_o;
  wire n603_o;
  wire n604_o;
  wire n605_o;
  wire [3:0] n606_o;
  wire n611_o;
  wire n612_o;
  wire n613_o;
  wire n614_o;
  wire n615_o;
  wire n616_o;
  wire n617_o;
  wire n618_o;
  wire n619_o;
  wire n620_o;
  wire n621_o;
  wire n622_o;
  wire n623_o;
  wire n624_o;
  wire n625_o;
  wire n626_o;
  wire n627_o;
  wire n628_o;
  wire n629_o;
  wire n630_o;
  wire n631_o;
  wire n632_o;
  wire n633_o;
  wire n634_o;
  wire n635_o;
  wire n636_o;
  wire n637_o;
  wire n638_o;
  wire [3:0] n639_o;
  wire n645_o;
  wire n646_o;
  wire n647_o;
  wire n648_o;
  wire n649_o;
  wire [3:0] n650_o;
  wire n657_o;
  wire n658_o;
  wire n659_o;
  wire n660_o;
  wire n661_o;
  wire [3:0] n662_o;
  wire n667_o;
  wire n668_o;
  wire n669_o;
  wire n670_o;
  wire n671_o;
  wire n672_o;
  wire n673_o;
  wire n674_o;
  wire n675_o;
  wire [3:0] n676_o;
  wire n682_o;
  wire n683_o;
  wire n684_o;
  wire n685_o;
  wire n686_o;
  wire [3:0] n687_o;
  wire n693_o;
  wire n694_o;
  wire n695_o;
  wire n696_o;
  wire n697_o;
  wire [3:0] n698_o;
  wire n704_o;
  wire n705_o;
  wire n706_o;
  wire n707_o;
  wire n708_o;
  wire [3:0] n709_o;
  wire [5:0] fsrom_block_fsroma;
  wire n717_o;
  wire n719_o;
  wire n721_o;
  wire n722_o;
  wire [4:0] n723_o;
  wire n724_o;
  wire n725_o;
  wire n726_o;
  wire [5:0] n727_o;
  wire n728_o;
  wire [3:0] n734_o;
  wire [1:0] n735_o;
  wire [5:0] n736_o;
  wire [5:0] n737_o;
  wire n740_o;
  wire n741_o;
  wire n742_o;
  wire n743_o;
  wire n744_o;
  wire n745_o;
  wire n746_o;
  wire n747_o;
  wire n748_o;
  wire n749_o;
  wire n750_o;
  wire n751_o;
  wire n752_o;
  wire n753_o;
  wire n754_o;
  wire n755_o;
  wire n756_o;
  wire n757_o;
  wire n758_o;
  wire n759_o;
  wire n760_o;
  wire n761_o;
  wire n762_o;
  wire n763_o;
  wire n764_o;
  wire n765_o;
  wire n766_o;
  wire n767_o;
  wire n768_o;
  wire n769_o;
  wire n770_o;
  wire n771_o;
  wire n772_o;
  wire n773_o;
  wire n774_o;
  wire n775_o;
  wire [5:0] fsrom_block_rom_block_na;
  wire [2:0] fsrom_block_rom_block_ndq;
  wire [17:0] fsrom_block_rom_block_wl;
  wire [5:0] n776_o;
  wire [2:0] n777_o;
  wire [2:0] n778_o;
  wire n779_o;
  wire n780_o;
  wire [1:0] n781_o;
  wire n782_o;
  wire [2:0] n783_o;
  wire n784_o;
  wire [3:0] n785_o;
  wire n786_o;
  wire [4:0] n787_o;
  wire n788_o;
  wire [5:0] n789_o;
  wire n790_o;
  wire [6:0] n791_o;
  wire n792_o;
  wire [7:0] n793_o;
  wire n794_o;
  wire [8:0] n795_o;
  wire n796_o;
  wire [9:0] n797_o;
  wire n798_o;
  wire [10:0] n799_o;
  wire n800_o;
  wire [11:0] n801_o;
  wire n802_o;
  wire [12:0] n803_o;
  wire n804_o;
  wire [13:0] n805_o;
  wire n806_o;
  wire [14:0] n807_o;
  wire n808_o;
  wire [15:0] n809_o;
  wire n810_o;
  wire [16:0] n811_o;
  wire n812_o;
  wire [17:0] n813_o;
  wire n820_o;
  wire n822_o;
  wire n824_o;
  wire n826_o;
  wire n828_o;
  wire n829_o;
  wire n830_o;
  wire n832_o;
  wire n833_o;
  wire n834_o;
  wire n836_o;
  wire n837_o;
  wire n838_o;
  wire n840_o;
  wire n841_o;
  wire n842_o;
  wire n844_o;
  wire n845_o;
  wire n846_o;
  wire n848_o;
  wire n849_o;
  wire n850_o;
  wire n852_o;
  wire n853_o;
  wire n854_o;
  wire n856_o;
  wire n857_o;
  wire n858_o;
  wire n860_o;
  wire n861_o;
  wire n862_o;
  wire n864_o;
  wire n865_o;
  wire n866_o;
  wire n868_o;
  wire n869_o;
  wire n870_o;
  wire n872_o;
  wire n873_o;
  wire n874_o;
  wire n876_o;
  wire n877_o;
  wire n878_o;
  wire n880_o;
  wire n881_o;
  wire n882_o;
  wire n884_o;
  wire n885_o;
  wire n886_o;
  wire n888_o;
  wire n889_o;
  wire n890_o;
  wire n892_o;
  wire n893_o;
  wire n894_o;
  wire n901_o;
  wire n903_o;
  wire n905_o;
  wire n907_o;
  wire n909_o;
  wire n910_o;
  wire n911_o;
  wire n913_o;
  wire n914_o;
  wire n915_o;
  wire n917_o;
  wire n918_o;
  wire n919_o;
  wire n921_o;
  wire n922_o;
  wire n923_o;
  wire n925_o;
  wire n926_o;
  wire n927_o;
  wire n929_o;
  wire n930_o;
  wire n931_o;
  wire n933_o;
  wire n934_o;
  wire n935_o;
  wire n937_o;
  wire n938_o;
  wire n939_o;
  wire n941_o;
  wire n942_o;
  wire n943_o;
  wire n945_o;
  wire n946_o;
  wire n947_o;
  wire n949_o;
  wire n950_o;
  wire n951_o;
  wire n953_o;
  wire n954_o;
  wire n955_o;
  wire n957_o;
  wire n958_o;
  wire n959_o;
  wire n961_o;
  wire n962_o;
  wire n963_o;
  wire n965_o;
  wire n966_o;
  wire n967_o;
  wire n969_o;
  wire n970_o;
  wire n971_o;
  wire n973_o;
  wire n974_o;
  wire n975_o;
  wire n982_o;
  wire n984_o;
  wire n986_o;
  wire n988_o;
  wire n990_o;
  wire n991_o;
  wire n992_o;
  wire n994_o;
  wire n995_o;
  wire n996_o;
  wire n998_o;
  wire n999_o;
  wire n1000_o;
  wire n1002_o;
  wire n1003_o;
  wire n1004_o;
  wire n1006_o;
  wire n1007_o;
  wire n1008_o;
  wire n1010_o;
  wire n1011_o;
  wire n1012_o;
  wire n1014_o;
  wire n1015_o;
  wire n1016_o;
  wire n1018_o;
  wire n1019_o;
  wire n1020_o;
  wire n1022_o;
  wire n1023_o;
  wire n1024_o;
  wire n1026_o;
  wire n1027_o;
  wire n1028_o;
  wire n1030_o;
  wire n1031_o;
  wire n1032_o;
  wire n1034_o;
  wire n1035_o;
  wire n1036_o;
  wire n1038_o;
  wire n1039_o;
  wire n1040_o;
  wire n1042_o;
  wire n1043_o;
  wire n1044_o;
  wire n1046_o;
  wire n1047_o;
  wire n1048_o;
  wire n1050_o;
  wire n1051_o;
  wire n1052_o;
  wire n1054_o;
  wire n1055_o;
  wire n1056_o;
  wire n1063_o;
  wire n1065_o;
  wire n1067_o;
  wire n1069_o;
  wire n1071_o;
  wire n1072_o;
  wire n1073_o;
  wire n1075_o;
  wire n1076_o;
  wire n1077_o;
  wire n1079_o;
  wire n1080_o;
  wire n1081_o;
  wire n1083_o;
  wire n1084_o;
  wire n1085_o;
  wire n1087_o;
  wire n1088_o;
  wire n1089_o;
  wire n1091_o;
  wire n1092_o;
  wire n1093_o;
  wire n1095_o;
  wire n1096_o;
  wire n1097_o;
  wire n1099_o;
  wire n1100_o;
  wire n1101_o;
  wire n1103_o;
  wire n1104_o;
  wire n1105_o;
  wire n1107_o;
  wire n1108_o;
  wire n1109_o;
  wire n1111_o;
  wire n1112_o;
  wire n1113_o;
  wire n1115_o;
  wire n1116_o;
  wire n1117_o;
  wire n1119_o;
  wire n1120_o;
  wire n1121_o;
  wire n1123_o;
  wire n1124_o;
  wire n1125_o;
  wire n1127_o;
  wire n1128_o;
  wire n1129_o;
  wire n1131_o;
  wire n1132_o;
  wire n1133_o;
  wire n1135_o;
  wire n1136_o;
  wire n1137_o;
  wire n1144_o;
  wire n1146_o;
  wire n1148_o;
  wire n1150_o;
  wire n1152_o;
  wire n1153_o;
  wire n1154_o;
  wire n1156_o;
  wire n1157_o;
  wire n1158_o;
  wire n1160_o;
  wire n1161_o;
  wire n1162_o;
  wire n1164_o;
  wire n1165_o;
  wire n1166_o;
  wire n1168_o;
  wire n1169_o;
  wire n1170_o;
  wire n1172_o;
  wire n1173_o;
  wire n1174_o;
  wire n1176_o;
  wire n1177_o;
  wire n1178_o;
  wire n1180_o;
  wire n1181_o;
  wire n1182_o;
  wire n1184_o;
  wire n1185_o;
  wire n1186_o;
  wire n1188_o;
  wire n1189_o;
  wire n1190_o;
  wire n1192_o;
  wire n1193_o;
  wire n1194_o;
  wire n1196_o;
  wire n1197_o;
  wire n1198_o;
  wire n1200_o;
  wire n1201_o;
  wire n1202_o;
  wire n1204_o;
  wire n1205_o;
  wire n1206_o;
  wire n1208_o;
  wire n1209_o;
  wire n1210_o;
  wire n1212_o;
  wire n1213_o;
  wire n1214_o;
  wire n1216_o;
  wire n1217_o;
  wire n1218_o;
  wire n1225_o;
  wire n1227_o;
  wire n1229_o;
  wire n1231_o;
  wire n1233_o;
  wire n1234_o;
  wire n1235_o;
  wire n1237_o;
  wire n1238_o;
  wire n1239_o;
  wire n1241_o;
  wire n1242_o;
  wire n1243_o;
  wire n1245_o;
  wire n1246_o;
  wire n1247_o;
  wire n1249_o;
  wire n1250_o;
  wire n1251_o;
  wire n1253_o;
  wire n1254_o;
  wire n1255_o;
  wire n1257_o;
  wire n1258_o;
  wire n1259_o;
  wire n1261_o;
  wire n1262_o;
  wire n1263_o;
  wire n1265_o;
  wire n1266_o;
  wire n1267_o;
  wire n1269_o;
  wire n1270_o;
  wire n1271_o;
  wire n1273_o;
  wire n1274_o;
  wire n1275_o;
  wire n1277_o;
  wire n1278_o;
  wire n1279_o;
  wire n1281_o;
  wire n1282_o;
  wire n1283_o;
  wire n1285_o;
  wire n1286_o;
  wire n1287_o;
  wire n1289_o;
  wire n1290_o;
  wire n1291_o;
  wire n1293_o;
  wire n1294_o;
  wire n1295_o;
  wire n1297_o;
  wire n1298_o;
  wire n1299_o;
  wire n1306_o;
  wire n1308_o;
  wire n1310_o;
  wire n1312_o;
  wire n1314_o;
  wire n1315_o;
  wire n1316_o;
  wire n1318_o;
  wire n1319_o;
  wire n1320_o;
  wire n1322_o;
  wire n1323_o;
  wire n1324_o;
  wire n1326_o;
  wire n1327_o;
  wire n1328_o;
  wire n1330_o;
  wire n1331_o;
  wire n1332_o;
  wire n1334_o;
  wire n1335_o;
  wire n1336_o;
  wire n1338_o;
  wire n1339_o;
  wire n1340_o;
  wire n1342_o;
  wire n1343_o;
  wire n1344_o;
  wire n1346_o;
  wire n1347_o;
  wire n1348_o;
  wire n1350_o;
  wire n1351_o;
  wire n1352_o;
  wire n1354_o;
  wire n1355_o;
  wire n1356_o;
  wire n1358_o;
  wire n1359_o;
  wire n1360_o;
  wire n1362_o;
  wire n1363_o;
  wire n1364_o;
  wire n1366_o;
  wire n1367_o;
  wire n1368_o;
  wire n1370_o;
  wire n1371_o;
  wire n1372_o;
  wire n1374_o;
  wire n1375_o;
  wire n1376_o;
  wire n1378_o;
  wire n1379_o;
  wire n1380_o;
  wire n1387_o;
  wire n1389_o;
  wire n1391_o;
  wire n1393_o;
  wire n1395_o;
  wire n1396_o;
  wire n1397_o;
  wire n1399_o;
  wire n1400_o;
  wire n1401_o;
  wire n1403_o;
  wire n1404_o;
  wire n1405_o;
  wire n1407_o;
  wire n1408_o;
  wire n1409_o;
  wire n1411_o;
  wire n1412_o;
  wire n1413_o;
  wire n1415_o;
  wire n1416_o;
  wire n1417_o;
  wire n1419_o;
  wire n1420_o;
  wire n1421_o;
  wire n1423_o;
  wire n1424_o;
  wire n1425_o;
  wire n1427_o;
  wire n1428_o;
  wire n1429_o;
  wire n1431_o;
  wire n1432_o;
  wire n1433_o;
  wire n1435_o;
  wire n1436_o;
  wire n1437_o;
  wire n1439_o;
  wire n1440_o;
  wire n1441_o;
  wire n1443_o;
  wire n1444_o;
  wire n1445_o;
  wire n1447_o;
  wire n1448_o;
  wire n1449_o;
  wire n1451_o;
  wire n1452_o;
  wire n1453_o;
  wire n1455_o;
  wire n1456_o;
  wire n1457_o;
  wire n1459_o;
  wire n1460_o;
  wire n1461_o;
  wire n1468_o;
  wire n1470_o;
  wire n1472_o;
  wire n1474_o;
  wire n1476_o;
  wire n1477_o;
  wire n1478_o;
  wire n1480_o;
  wire n1481_o;
  wire n1482_o;
  wire n1484_o;
  wire n1485_o;
  wire n1486_o;
  wire n1488_o;
  wire n1489_o;
  wire n1490_o;
  wire n1492_o;
  wire n1493_o;
  wire n1494_o;
  wire n1496_o;
  wire n1497_o;
  wire n1498_o;
  wire n1500_o;
  wire n1501_o;
  wire n1502_o;
  wire n1504_o;
  wire n1505_o;
  wire n1506_o;
  wire n1508_o;
  wire n1509_o;
  wire n1510_o;
  wire n1512_o;
  wire n1513_o;
  wire n1514_o;
  wire n1516_o;
  wire n1517_o;
  wire n1518_o;
  wire n1520_o;
  wire n1521_o;
  wire n1522_o;
  wire n1524_o;
  wire n1525_o;
  wire n1526_o;
  wire n1528_o;
  wire n1529_o;
  wire n1530_o;
  wire n1532_o;
  wire n1533_o;
  wire n1534_o;
  wire n1536_o;
  wire n1537_o;
  wire n1538_o;
  wire n1540_o;
  wire n1541_o;
  wire n1542_o;
  wire n1549_o;
  wire n1551_o;
  wire n1553_o;
  wire n1555_o;
  wire n1557_o;
  wire n1558_o;
  wire n1559_o;
  wire n1561_o;
  wire n1562_o;
  wire n1563_o;
  wire n1565_o;
  wire n1566_o;
  wire n1567_o;
  wire n1569_o;
  wire n1570_o;
  wire n1571_o;
  wire n1573_o;
  wire n1574_o;
  wire n1575_o;
  wire n1577_o;
  wire n1578_o;
  wire n1579_o;
  wire n1581_o;
  wire n1582_o;
  wire n1583_o;
  wire n1585_o;
  wire n1586_o;
  wire n1587_o;
  wire n1589_o;
  wire n1590_o;
  wire n1591_o;
  wire n1593_o;
  wire n1594_o;
  wire n1595_o;
  wire n1597_o;
  wire n1598_o;
  wire n1599_o;
  wire n1601_o;
  wire n1602_o;
  wire n1603_o;
  wire n1605_o;
  wire n1606_o;
  wire n1607_o;
  wire n1609_o;
  wire n1610_o;
  wire n1611_o;
  wire n1613_o;
  wire n1614_o;
  wire n1615_o;
  wire n1617_o;
  wire n1618_o;
  wire n1619_o;
  wire n1621_o;
  wire n1622_o;
  wire n1623_o;
  wire n1630_o;
  wire n1632_o;
  wire n1634_o;
  wire n1636_o;
  wire n1638_o;
  wire n1639_o;
  wire n1640_o;
  wire n1642_o;
  wire n1643_o;
  wire n1644_o;
  wire n1646_o;
  wire n1647_o;
  wire n1648_o;
  wire n1650_o;
  wire n1651_o;
  wire n1652_o;
  wire n1654_o;
  wire n1655_o;
  wire n1656_o;
  wire n1658_o;
  wire n1659_o;
  wire n1660_o;
  wire n1662_o;
  wire n1663_o;
  wire n1664_o;
  wire n1666_o;
  wire n1667_o;
  wire n1668_o;
  wire n1670_o;
  wire n1671_o;
  wire n1672_o;
  wire n1674_o;
  wire n1675_o;
  wire n1676_o;
  wire n1678_o;
  wire n1679_o;
  wire n1680_o;
  wire n1682_o;
  wire n1683_o;
  wire n1684_o;
  wire n1686_o;
  wire n1687_o;
  wire n1688_o;
  wire n1690_o;
  wire n1691_o;
  wire n1692_o;
  wire n1694_o;
  wire n1695_o;
  wire n1696_o;
  wire n1698_o;
  wire n1699_o;
  wire n1700_o;
  wire n1702_o;
  wire n1703_o;
  wire n1704_o;
  wire n1711_o;
  wire n1713_o;
  wire n1715_o;
  wire n1717_o;
  wire n1719_o;
  wire n1720_o;
  wire n1721_o;
  wire n1723_o;
  wire n1724_o;
  wire n1725_o;
  wire n1727_o;
  wire n1728_o;
  wire n1729_o;
  wire n1731_o;
  wire n1732_o;
  wire n1733_o;
  wire n1735_o;
  wire n1736_o;
  wire n1737_o;
  wire n1739_o;
  wire n1740_o;
  wire n1741_o;
  wire n1743_o;
  wire n1744_o;
  wire n1745_o;
  wire n1747_o;
  wire n1748_o;
  wire n1749_o;
  wire n1751_o;
  wire n1752_o;
  wire n1753_o;
  wire n1755_o;
  wire n1756_o;
  wire n1757_o;
  wire n1759_o;
  wire n1760_o;
  wire n1761_o;
  wire n1763_o;
  wire n1764_o;
  wire n1765_o;
  wire n1767_o;
  wire n1768_o;
  wire n1769_o;
  wire n1771_o;
  wire n1772_o;
  wire n1773_o;
  wire n1775_o;
  wire n1776_o;
  wire n1777_o;
  wire n1779_o;
  wire n1780_o;
  wire n1781_o;
  wire n1783_o;
  wire n1784_o;
  wire n1785_o;
  wire n1792_o;
  wire n1794_o;
  wire n1796_o;
  wire n1798_o;
  wire n1800_o;
  wire n1801_o;
  wire n1802_o;
  wire n1804_o;
  wire n1805_o;
  wire n1806_o;
  wire n1808_o;
  wire n1809_o;
  wire n1810_o;
  wire n1812_o;
  wire n1813_o;
  wire n1814_o;
  wire n1816_o;
  wire n1817_o;
  wire n1818_o;
  wire n1820_o;
  wire n1821_o;
  wire n1822_o;
  wire n1824_o;
  wire n1825_o;
  wire n1826_o;
  wire n1828_o;
  wire n1829_o;
  wire n1830_o;
  wire n1832_o;
  wire n1833_o;
  wire n1834_o;
  wire n1836_o;
  wire n1837_o;
  wire n1838_o;
  wire n1840_o;
  wire n1841_o;
  wire n1842_o;
  wire n1844_o;
  wire n1845_o;
  wire n1846_o;
  wire n1848_o;
  wire n1849_o;
  wire n1850_o;
  wire n1852_o;
  wire n1853_o;
  wire n1854_o;
  wire n1856_o;
  wire n1857_o;
  wire n1858_o;
  wire n1860_o;
  wire n1861_o;
  wire n1862_o;
  wire n1864_o;
  wire n1865_o;
  wire n1866_o;
  wire n1873_o;
  wire n1875_o;
  wire n1877_o;
  wire n1879_o;
  wire n1881_o;
  wire n1882_o;
  wire n1883_o;
  wire n1885_o;
  wire n1886_o;
  wire n1887_o;
  wire n1889_o;
  wire n1890_o;
  wire n1891_o;
  wire n1893_o;
  wire n1894_o;
  wire n1895_o;
  wire n1897_o;
  wire n1898_o;
  wire n1899_o;
  wire n1901_o;
  wire n1902_o;
  wire n1903_o;
  wire n1905_o;
  wire n1906_o;
  wire n1907_o;
  wire n1909_o;
  wire n1910_o;
  wire n1911_o;
  wire n1913_o;
  wire n1914_o;
  wire n1915_o;
  wire n1917_o;
  wire n1918_o;
  wire n1919_o;
  wire n1921_o;
  wire n1922_o;
  wire n1923_o;
  wire n1925_o;
  wire n1926_o;
  wire n1927_o;
  wire n1929_o;
  wire n1930_o;
  wire n1931_o;
  wire n1933_o;
  wire n1934_o;
  wire n1935_o;
  wire n1937_o;
  wire n1938_o;
  wire n1939_o;
  wire n1941_o;
  wire n1942_o;
  wire n1943_o;
  wire n1945_o;
  wire n1946_o;
  wire n1947_o;
  wire [3:0] n1948_o;
  wire [3:0] n1949_o;
  wire [3:0] n1950_o;
  wire [1:0] n1951_o;
  wire [13:0] n1952_o;
  wire [5:0] n1954_o;
  wire n1960_o;
  wire n1962_o;
  wire n1964_o;
  wire n1965_o;
  wire n1966_o;
  wire n1967_o;
  wire n1968_o;
  wire n1969_o;
  wire n1970_o;
  wire n1971_o;
  wire n1972_o;
  wire n1973_o;
  wire n1974_o;
  wire [5:0] n1976_o;
  wire n1982_o;
  wire n1984_o;
  wire n1986_o;
  wire n1987_o;
  wire n1988_o;
  wire n1989_o;
  wire n1990_o;
  wire n1991_o;
  wire n1992_o;
  wire n1993_o;
  wire n1994_o;
  wire n1995_o;
  wire n1996_o;
  wire [5:0] n1997_o;
  reg [5:0] n1998_q;
  wire [4:0] seqrom_block_gseqroma;
  wire seqrom_block_agen_block_ncen3;
  reg [4:0] seqrom_block_agen_block_seqroma;
  wire n2005_o;
  wire n2006_o;
  wire n2012_o;
  wire n2013_o;
  wire n2014_o;
  wire n2015_o;
  wire n2016_o;
  wire n2017_o;
  wire n2018_o;
  wire n2019_o;
  wire n2020_o;
  wire [3:0] n2021_o;
  wire n2022_o;
  wire n2023_o;
  wire n2024_o;
  wire n2032_o;
  wire n2034_o;
  wire n2036_o;
  wire n2037_o;
  wire n2038_o;
  wire n2039_o;
  wire n2040_o;
  wire n2041_o;
  wire n2042_o;
  wire n2043_o;
  wire n2044_o;
  wire n2045_o;
  wire n2046_o;
  wire n2047_o;
  wire n2048_o;
  wire n2049_o;
  wire n2050_o;
  wire n2051_o;
  wire [3:0] n2052_o;
  wire [3:0] n2053_o;
  wire [3:0] n2054_o;
  wire n2055_o;
  wire [3:0] n2057_o;
  wire n2058_o;
  wire [4:0] n2060_o;
  wire n2063_o;
  wire [3:0] n2064_o;
  wire n2065_o;
  wire n2066_o;
  wire [4:0] n2067_o;
  wire n2068_o;
  wire [4:0] n2069_o;
  reg [4:0] n2070_q;
  wire [4:0] seqrom_block_rom_block_na;
  wire [4:0] seqrom_block_rom_block_ny;
  wire [11:0] seqrom_block_rom_block_xwl;
  wire [35:0] seqrom_block_rom_block_ywl;
  wire [4:0] n2071_o;
  wire n2072_o;
  wire n2073_o;
  wire [1:0] n2074_o;
  wire n2075_o;
  wire [2:0] n2076_o;
  wire n2077_o;
  wire [3:0] n2078_o;
  wire n2079_o;
  wire [4:0] n2080_o;
  wire n2081_o;
  wire [5:0] n2082_o;
  wire n2083_o;
  wire [6:0] n2084_o;
  wire n2085_o;
  wire [7:0] n2086_o;
  wire n2087_o;
  wire [8:0] n2088_o;
  wire n2089_o;
  wire [9:0] n2090_o;
  wire n2091_o;
  wire [10:0] n2092_o;
  wire n2093_o;
  wire [11:0] n2094_o;
  wire n2101_o;
  wire n2103_o;
  wire n2105_o;
  wire n2107_o;
  wire n2109_o;
  wire n2110_o;
  wire n2111_o;
  wire n2113_o;
  wire n2114_o;
  wire n2115_o;
  wire n2117_o;
  wire n2118_o;
  wire n2119_o;
  wire n2121_o;
  wire n2122_o;
  wire n2123_o;
  wire n2125_o;
  wire n2126_o;
  wire n2127_o;
  wire n2129_o;
  wire n2130_o;
  wire n2131_o;
  wire n2133_o;
  wire n2134_o;
  wire n2135_o;
  wire n2137_o;
  wire n2138_o;
  wire n2139_o;
  wire n2141_o;
  wire n2142_o;
  wire n2143_o;
  wire n2145_o;
  wire n2146_o;
  wire n2147_o;
  wire n2149_o;
  wire n2150_o;
  wire n2151_o;
  wire n2158_o;
  wire n2160_o;
  wire n2162_o;
  wire n2164_o;
  wire n2166_o;
  wire n2167_o;
  wire n2168_o;
  wire n2170_o;
  wire n2171_o;
  wire n2172_o;
  wire n2174_o;
  wire n2175_o;
  wire n2176_o;
  wire n2178_o;
  wire n2179_o;
  wire n2180_o;
  wire n2182_o;
  wire n2183_o;
  wire n2184_o;
  wire n2186_o;
  wire n2187_o;
  wire n2188_o;
  wire n2190_o;
  wire n2191_o;
  wire n2192_o;
  wire n2194_o;
  wire n2195_o;
  wire n2196_o;
  wire n2198_o;
  wire n2199_o;
  wire n2200_o;
  wire n2202_o;
  wire n2203_o;
  wire n2204_o;
  wire n2206_o;
  wire n2207_o;
  wire n2208_o;
  wire n2215_o;
  wire n2217_o;
  wire n2219_o;
  wire n2221_o;
  wire n2223_o;
  wire n2224_o;
  wire n2225_o;
  wire n2227_o;
  wire n2228_o;
  wire n2229_o;
  wire n2231_o;
  wire n2232_o;
  wire n2233_o;
  wire n2235_o;
  wire n2236_o;
  wire n2237_o;
  wire n2239_o;
  wire n2240_o;
  wire n2241_o;
  wire n2243_o;
  wire n2244_o;
  wire n2245_o;
  wire n2247_o;
  wire n2248_o;
  wire n2249_o;
  wire n2251_o;
  wire n2252_o;
  wire n2253_o;
  wire n2255_o;
  wire n2256_o;
  wire n2257_o;
  wire n2259_o;
  wire n2260_o;
  wire n2261_o;
  wire n2263_o;
  wire n2264_o;
  wire n2265_o;
  wire n2272_o;
  wire n2274_o;
  wire n2276_o;
  wire n2278_o;
  wire n2280_o;
  wire n2281_o;
  wire n2282_o;
  wire n2284_o;
  wire n2285_o;
  wire n2286_o;
  wire n2288_o;
  wire n2289_o;
  wire n2290_o;
  wire n2292_o;
  wire n2293_o;
  wire n2294_o;
  wire n2296_o;
  wire n2297_o;
  wire n2298_o;
  wire n2300_o;
  wire n2301_o;
  wire n2302_o;
  wire n2304_o;
  wire n2305_o;
  wire n2306_o;
  wire n2308_o;
  wire n2309_o;
  wire n2310_o;
  wire n2312_o;
  wire n2313_o;
  wire n2314_o;
  wire n2316_o;
  wire n2317_o;
  wire n2318_o;
  wire n2320_o;
  wire n2321_o;
  wire n2322_o;
  wire n2329_o;
  wire n2331_o;
  wire n2333_o;
  wire n2335_o;
  wire n2337_o;
  wire n2338_o;
  wire n2339_o;
  wire n2341_o;
  wire n2342_o;
  wire n2343_o;
  wire n2345_o;
  wire n2346_o;
  wire n2347_o;
  wire n2349_o;
  wire n2350_o;
  wire n2351_o;
  wire n2353_o;
  wire n2354_o;
  wire n2355_o;
  wire n2357_o;
  wire n2358_o;
  wire n2359_o;
  wire n2361_o;
  wire n2362_o;
  wire n2363_o;
  wire n2365_o;
  wire n2366_o;
  wire n2367_o;
  wire n2369_o;
  wire n2370_o;
  wire n2371_o;
  wire n2373_o;
  wire n2374_o;
  wire n2375_o;
  wire n2377_o;
  wire n2378_o;
  wire n2379_o;
  wire n2386_o;
  wire n2388_o;
  wire n2390_o;
  wire n2392_o;
  wire n2394_o;
  wire n2395_o;
  wire n2396_o;
  wire n2398_o;
  wire n2399_o;
  wire n2400_o;
  wire n2402_o;
  wire n2403_o;
  wire n2404_o;
  wire n2406_o;
  wire n2407_o;
  wire n2408_o;
  wire n2410_o;
  wire n2411_o;
  wire n2412_o;
  wire n2414_o;
  wire n2415_o;
  wire n2416_o;
  wire n2418_o;
  wire n2419_o;
  wire n2420_o;
  wire n2422_o;
  wire n2423_o;
  wire n2424_o;
  wire n2426_o;
  wire n2427_o;
  wire n2428_o;
  wire n2430_o;
  wire n2431_o;
  wire n2432_o;
  wire n2434_o;
  wire n2435_o;
  wire n2436_o;
  wire n2443_o;
  wire n2445_o;
  wire n2447_o;
  wire n2449_o;
  wire n2451_o;
  wire n2452_o;
  wire n2453_o;
  wire n2455_o;
  wire n2456_o;
  wire n2457_o;
  wire n2459_o;
  wire n2460_o;
  wire n2461_o;
  wire n2463_o;
  wire n2464_o;
  wire n2465_o;
  wire n2467_o;
  wire n2468_o;
  wire n2469_o;
  wire n2471_o;
  wire n2472_o;
  wire n2473_o;
  wire n2475_o;
  wire n2476_o;
  wire n2477_o;
  wire n2479_o;
  wire n2480_o;
  wire n2481_o;
  wire n2483_o;
  wire n2484_o;
  wire n2485_o;
  wire n2487_o;
  wire n2488_o;
  wire n2489_o;
  wire n2491_o;
  wire n2492_o;
  wire n2493_o;
  wire n2500_o;
  wire n2502_o;
  wire n2504_o;
  wire n2506_o;
  wire n2508_o;
  wire n2509_o;
  wire n2510_o;
  wire n2512_o;
  wire n2513_o;
  wire n2514_o;
  wire n2516_o;
  wire n2517_o;
  wire n2518_o;
  wire n2520_o;
  wire n2521_o;
  wire n2522_o;
  wire n2524_o;
  wire n2525_o;
  wire n2526_o;
  wire n2528_o;
  wire n2529_o;
  wire n2530_o;
  wire n2532_o;
  wire n2533_o;
  wire n2534_o;
  wire n2536_o;
  wire n2537_o;
  wire n2538_o;
  wire n2540_o;
  wire n2541_o;
  wire n2542_o;
  wire n2544_o;
  wire n2545_o;
  wire n2546_o;
  wire n2548_o;
  wire n2549_o;
  wire n2550_o;
  wire n2557_o;
  wire n2559_o;
  wire n2561_o;
  wire n2563_o;
  wire n2565_o;
  wire n2566_o;
  wire n2567_o;
  wire n2569_o;
  wire n2570_o;
  wire n2571_o;
  wire n2573_o;
  wire n2574_o;
  wire n2575_o;
  wire n2577_o;
  wire n2578_o;
  wire n2579_o;
  wire n2581_o;
  wire n2582_o;
  wire n2583_o;
  wire n2585_o;
  wire n2586_o;
  wire n2587_o;
  wire n2589_o;
  wire n2590_o;
  wire n2591_o;
  wire n2593_o;
  wire n2594_o;
  wire n2595_o;
  wire n2597_o;
  wire n2598_o;
  wire n2599_o;
  wire n2601_o;
  wire n2602_o;
  wire n2603_o;
  wire n2605_o;
  wire n2606_o;
  wire n2607_o;
  wire n2614_o;
  wire n2616_o;
  wire n2618_o;
  wire n2620_o;
  wire n2622_o;
  wire n2623_o;
  wire n2624_o;
  wire n2626_o;
  wire n2627_o;
  wire n2628_o;
  wire n2630_o;
  wire n2631_o;
  wire n2632_o;
  wire n2634_o;
  wire n2635_o;
  wire n2636_o;
  wire n2638_o;
  wire n2639_o;
  wire n2640_o;
  wire n2642_o;
  wire n2643_o;
  wire n2644_o;
  wire n2646_o;
  wire n2647_o;
  wire n2648_o;
  wire n2650_o;
  wire n2651_o;
  wire n2652_o;
  wire n2654_o;
  wire n2655_o;
  wire n2656_o;
  wire n2658_o;
  wire n2659_o;
  wire n2660_o;
  wire n2662_o;
  wire n2663_o;
  wire n2664_o;
  wire n2671_o;
  wire n2673_o;
  wire n2675_o;
  wire n2677_o;
  wire n2679_o;
  wire n2680_o;
  wire n2681_o;
  wire n2683_o;
  wire n2684_o;
  wire n2685_o;
  wire n2687_o;
  wire n2688_o;
  wire n2689_o;
  wire n2691_o;
  wire n2692_o;
  wire n2693_o;
  wire n2695_o;
  wire n2696_o;
  wire n2697_o;
  wire n2699_o;
  wire n2700_o;
  wire n2701_o;
  wire n2703_o;
  wire n2704_o;
  wire n2705_o;
  wire n2707_o;
  wire n2708_o;
  wire n2709_o;
  wire n2711_o;
  wire n2712_o;
  wire n2713_o;
  wire n2715_o;
  wire n2716_o;
  wire n2717_o;
  wire n2719_o;
  wire n2720_o;
  wire n2721_o;
  wire n2728_o;
  wire n2730_o;
  wire n2732_o;
  wire n2734_o;
  wire n2736_o;
  wire n2737_o;
  wire n2738_o;
  wire n2740_o;
  wire n2741_o;
  wire n2742_o;
  wire n2744_o;
  wire n2745_o;
  wire n2746_o;
  wire n2748_o;
  wire n2749_o;
  wire n2750_o;
  wire n2752_o;
  wire n2753_o;
  wire n2754_o;
  wire n2756_o;
  wire n2757_o;
  wire n2758_o;
  wire n2760_o;
  wire n2761_o;
  wire n2762_o;
  wire n2764_o;
  wire n2765_o;
  wire n2766_o;
  wire n2768_o;
  wire n2769_o;
  wire n2770_o;
  wire n2772_o;
  wire n2773_o;
  wire n2774_o;
  wire n2776_o;
  wire n2777_o;
  wire n2778_o;
  wire n2785_o;
  wire n2787_o;
  wire n2789_o;
  wire n2791_o;
  wire n2793_o;
  wire n2794_o;
  wire n2795_o;
  wire n2797_o;
  wire n2798_o;
  wire n2799_o;
  wire n2801_o;
  wire n2802_o;
  wire n2803_o;
  wire n2805_o;
  wire n2806_o;
  wire n2807_o;
  wire n2809_o;
  wire n2810_o;
  wire n2811_o;
  wire n2813_o;
  wire n2814_o;
  wire n2815_o;
  wire n2817_o;
  wire n2818_o;
  wire n2819_o;
  wire n2821_o;
  wire n2822_o;
  wire n2823_o;
  wire n2825_o;
  wire n2826_o;
  wire n2827_o;
  wire n2829_o;
  wire n2830_o;
  wire n2831_o;
  wire n2833_o;
  wire n2834_o;
  wire n2835_o;
  wire n2842_o;
  wire n2844_o;
  wire n2846_o;
  wire n2848_o;
  wire n2850_o;
  wire n2851_o;
  wire n2852_o;
  wire n2854_o;
  wire n2855_o;
  wire n2856_o;
  wire n2858_o;
  wire n2859_o;
  wire n2860_o;
  wire n2862_o;
  wire n2863_o;
  wire n2864_o;
  wire n2866_o;
  wire n2867_o;
  wire n2868_o;
  wire n2870_o;
  wire n2871_o;
  wire n2872_o;
  wire n2874_o;
  wire n2875_o;
  wire n2876_o;
  wire n2878_o;
  wire n2879_o;
  wire n2880_o;
  wire n2882_o;
  wire n2883_o;
  wire n2884_o;
  wire n2886_o;
  wire n2887_o;
  wire n2888_o;
  wire n2890_o;
  wire n2891_o;
  wire n2892_o;
  wire n2899_o;
  wire n2901_o;
  wire n2903_o;
  wire n2905_o;
  wire n2907_o;
  wire n2908_o;
  wire n2909_o;
  wire n2911_o;
  wire n2912_o;
  wire n2913_o;
  wire n2915_o;
  wire n2916_o;
  wire n2917_o;
  wire n2919_o;
  wire n2920_o;
  wire n2921_o;
  wire n2923_o;
  wire n2924_o;
  wire n2925_o;
  wire n2927_o;
  wire n2928_o;
  wire n2929_o;
  wire n2931_o;
  wire n2932_o;
  wire n2933_o;
  wire n2935_o;
  wire n2936_o;
  wire n2937_o;
  wire n2939_o;
  wire n2940_o;
  wire n2941_o;
  wire n2943_o;
  wire n2944_o;
  wire n2945_o;
  wire n2947_o;
  wire n2948_o;
  wire n2949_o;
  wire n2956_o;
  wire n2958_o;
  wire n2960_o;
  wire n2962_o;
  wire n2964_o;
  wire n2965_o;
  wire n2966_o;
  wire n2968_o;
  wire n2969_o;
  wire n2970_o;
  wire n2972_o;
  wire n2973_o;
  wire n2974_o;
  wire n2976_o;
  wire n2977_o;
  wire n2978_o;
  wire n2980_o;
  wire n2981_o;
  wire n2982_o;
  wire n2984_o;
  wire n2985_o;
  wire n2986_o;
  wire n2988_o;
  wire n2989_o;
  wire n2990_o;
  wire n2992_o;
  wire n2993_o;
  wire n2994_o;
  wire n2996_o;
  wire n2997_o;
  wire n2998_o;
  wire n3000_o;
  wire n3001_o;
  wire n3002_o;
  wire n3004_o;
  wire n3005_o;
  wire n3006_o;
  wire n3013_o;
  wire n3015_o;
  wire n3017_o;
  wire n3019_o;
  wire n3021_o;
  wire n3022_o;
  wire n3023_o;
  wire n3025_o;
  wire n3026_o;
  wire n3027_o;
  wire n3029_o;
  wire n3030_o;
  wire n3031_o;
  wire n3033_o;
  wire n3034_o;
  wire n3035_o;
  wire n3037_o;
  wire n3038_o;
  wire n3039_o;
  wire n3041_o;
  wire n3042_o;
  wire n3043_o;
  wire n3045_o;
  wire n3046_o;
  wire n3047_o;
  wire n3049_o;
  wire n3050_o;
  wire n3051_o;
  wire n3053_o;
  wire n3054_o;
  wire n3055_o;
  wire n3057_o;
  wire n3058_o;
  wire n3059_o;
  wire n3061_o;
  wire n3062_o;
  wire n3063_o;
  wire n3070_o;
  wire n3072_o;
  wire n3074_o;
  wire n3076_o;
  wire n3078_o;
  wire n3079_o;
  wire n3080_o;
  wire n3082_o;
  wire n3083_o;
  wire n3084_o;
  wire n3086_o;
  wire n3087_o;
  wire n3088_o;
  wire n3090_o;
  wire n3091_o;
  wire n3092_o;
  wire n3094_o;
  wire n3095_o;
  wire n3096_o;
  wire n3098_o;
  wire n3099_o;
  wire n3100_o;
  wire n3102_o;
  wire n3103_o;
  wire n3104_o;
  wire n3106_o;
  wire n3107_o;
  wire n3108_o;
  wire n3110_o;
  wire n3111_o;
  wire n3112_o;
  wire n3114_o;
  wire n3115_o;
  wire n3116_o;
  wire n3118_o;
  wire n3119_o;
  wire n3120_o;
  wire n3127_o;
  wire n3129_o;
  wire n3131_o;
  wire n3133_o;
  wire n3135_o;
  wire n3136_o;
  wire n3137_o;
  wire n3139_o;
  wire n3140_o;
  wire n3141_o;
  wire n3143_o;
  wire n3144_o;
  wire n3145_o;
  wire n3147_o;
  wire n3148_o;
  wire n3149_o;
  wire n3151_o;
  wire n3152_o;
  wire n3153_o;
  wire n3155_o;
  wire n3156_o;
  wire n3157_o;
  wire n3159_o;
  wire n3160_o;
  wire n3161_o;
  wire n3163_o;
  wire n3164_o;
  wire n3165_o;
  wire n3167_o;
  wire n3168_o;
  wire n3169_o;
  wire n3171_o;
  wire n3172_o;
  wire n3173_o;
  wire n3175_o;
  wire n3176_o;
  wire n3177_o;
  wire n3184_o;
  wire n3186_o;
  wire n3188_o;
  wire n3190_o;
  wire n3192_o;
  wire n3193_o;
  wire n3194_o;
  wire n3196_o;
  wire n3197_o;
  wire n3198_o;
  wire n3200_o;
  wire n3201_o;
  wire n3202_o;
  wire n3204_o;
  wire n3205_o;
  wire n3206_o;
  wire n3208_o;
  wire n3209_o;
  wire n3210_o;
  wire n3212_o;
  wire n3213_o;
  wire n3214_o;
  wire n3216_o;
  wire n3217_o;
  wire n3218_o;
  wire n3220_o;
  wire n3221_o;
  wire n3222_o;
  wire n3224_o;
  wire n3225_o;
  wire n3226_o;
  wire n3228_o;
  wire n3229_o;
  wire n3230_o;
  wire n3232_o;
  wire n3233_o;
  wire n3234_o;
  wire n3241_o;
  wire n3243_o;
  wire n3245_o;
  wire n3247_o;
  wire n3249_o;
  wire n3250_o;
  wire n3251_o;
  wire n3253_o;
  wire n3254_o;
  wire n3255_o;
  wire n3257_o;
  wire n3258_o;
  wire n3259_o;
  wire n3261_o;
  wire n3262_o;
  wire n3263_o;
  wire n3265_o;
  wire n3266_o;
  wire n3267_o;
  wire n3269_o;
  wire n3270_o;
  wire n3271_o;
  wire n3273_o;
  wire n3274_o;
  wire n3275_o;
  wire n3277_o;
  wire n3278_o;
  wire n3279_o;
  wire n3281_o;
  wire n3282_o;
  wire n3283_o;
  wire n3285_o;
  wire n3286_o;
  wire n3287_o;
  wire n3289_o;
  wire n3290_o;
  wire n3291_o;
  wire n3298_o;
  wire n3300_o;
  wire n3302_o;
  wire n3304_o;
  wire n3306_o;
  wire n3307_o;
  wire n3308_o;
  wire n3310_o;
  wire n3311_o;
  wire n3312_o;
  wire n3314_o;
  wire n3315_o;
  wire n3316_o;
  wire n3318_o;
  wire n3319_o;
  wire n3320_o;
  wire n3322_o;
  wire n3323_o;
  wire n3324_o;
  wire n3326_o;
  wire n3327_o;
  wire n3328_o;
  wire n3330_o;
  wire n3331_o;
  wire n3332_o;
  wire n3334_o;
  wire n3335_o;
  wire n3336_o;
  wire n3338_o;
  wire n3339_o;
  wire n3340_o;
  wire n3342_o;
  wire n3343_o;
  wire n3344_o;
  wire n3346_o;
  wire n3347_o;
  wire n3348_o;
  wire n3355_o;
  wire n3357_o;
  wire n3359_o;
  wire n3361_o;
  wire n3363_o;
  wire n3364_o;
  wire n3365_o;
  wire n3367_o;
  wire n3368_o;
  wire n3369_o;
  wire n3371_o;
  wire n3372_o;
  wire n3373_o;
  wire n3375_o;
  wire n3376_o;
  wire n3377_o;
  wire n3379_o;
  wire n3380_o;
  wire n3381_o;
  wire n3383_o;
  wire n3384_o;
  wire n3385_o;
  wire n3387_o;
  wire n3388_o;
  wire n3389_o;
  wire n3391_o;
  wire n3392_o;
  wire n3393_o;
  wire n3395_o;
  wire n3396_o;
  wire n3397_o;
  wire n3399_o;
  wire n3400_o;
  wire n3401_o;
  wire n3403_o;
  wire n3404_o;
  wire n3405_o;
  wire n3412_o;
  wire n3414_o;
  wire n3416_o;
  wire n3418_o;
  wire n3420_o;
  wire n3421_o;
  wire n3422_o;
  wire n3424_o;
  wire n3425_o;
  wire n3426_o;
  wire n3428_o;
  wire n3429_o;
  wire n3430_o;
  wire n3432_o;
  wire n3433_o;
  wire n3434_o;
  wire n3436_o;
  wire n3437_o;
  wire n3438_o;
  wire n3440_o;
  wire n3441_o;
  wire n3442_o;
  wire n3444_o;
  wire n3445_o;
  wire n3446_o;
  wire n3448_o;
  wire n3449_o;
  wire n3450_o;
  wire n3452_o;
  wire n3453_o;
  wire n3454_o;
  wire n3456_o;
  wire n3457_o;
  wire n3458_o;
  wire n3460_o;
  wire n3461_o;
  wire n3462_o;
  wire n3469_o;
  wire n3471_o;
  wire n3473_o;
  wire n3475_o;
  wire n3477_o;
  wire n3478_o;
  wire n3479_o;
  wire n3481_o;
  wire n3482_o;
  wire n3483_o;
  wire n3485_o;
  wire n3486_o;
  wire n3487_o;
  wire n3489_o;
  wire n3490_o;
  wire n3491_o;
  wire n3493_o;
  wire n3494_o;
  wire n3495_o;
  wire n3497_o;
  wire n3498_o;
  wire n3499_o;
  wire n3501_o;
  wire n3502_o;
  wire n3503_o;
  wire n3505_o;
  wire n3506_o;
  wire n3507_o;
  wire n3509_o;
  wire n3510_o;
  wire n3511_o;
  wire n3513_o;
  wire n3514_o;
  wire n3515_o;
  wire n3517_o;
  wire n3518_o;
  wire n3519_o;
  wire n3526_o;
  wire n3528_o;
  wire n3530_o;
  wire n3532_o;
  wire n3534_o;
  wire n3535_o;
  wire n3536_o;
  wire n3538_o;
  wire n3539_o;
  wire n3540_o;
  wire n3542_o;
  wire n3543_o;
  wire n3544_o;
  wire n3546_o;
  wire n3547_o;
  wire n3548_o;
  wire n3550_o;
  wire n3551_o;
  wire n3552_o;
  wire n3554_o;
  wire n3555_o;
  wire n3556_o;
  wire n3558_o;
  wire n3559_o;
  wire n3560_o;
  wire n3562_o;
  wire n3563_o;
  wire n3564_o;
  wire n3566_o;
  wire n3567_o;
  wire n3568_o;
  wire n3570_o;
  wire n3571_o;
  wire n3572_o;
  wire n3574_o;
  wire n3575_o;
  wire n3576_o;
  wire n3583_o;
  wire n3585_o;
  wire n3587_o;
  wire n3589_o;
  wire n3591_o;
  wire n3592_o;
  wire n3593_o;
  wire n3595_o;
  wire n3596_o;
  wire n3597_o;
  wire n3599_o;
  wire n3600_o;
  wire n3601_o;
  wire n3603_o;
  wire n3604_o;
  wire n3605_o;
  wire n3607_o;
  wire n3608_o;
  wire n3609_o;
  wire n3611_o;
  wire n3612_o;
  wire n3613_o;
  wire n3615_o;
  wire n3616_o;
  wire n3617_o;
  wire n3619_o;
  wire n3620_o;
  wire n3621_o;
  wire n3623_o;
  wire n3624_o;
  wire n3625_o;
  wire n3627_o;
  wire n3628_o;
  wire n3629_o;
  wire n3631_o;
  wire n3632_o;
  wire n3633_o;
  wire n3640_o;
  wire n3642_o;
  wire n3644_o;
  wire n3646_o;
  wire n3648_o;
  wire n3649_o;
  wire n3650_o;
  wire n3652_o;
  wire n3653_o;
  wire n3654_o;
  wire n3656_o;
  wire n3657_o;
  wire n3658_o;
  wire n3660_o;
  wire n3661_o;
  wire n3662_o;
  wire n3664_o;
  wire n3665_o;
  wire n3666_o;
  wire n3668_o;
  wire n3669_o;
  wire n3670_o;
  wire n3672_o;
  wire n3673_o;
  wire n3674_o;
  wire n3676_o;
  wire n3677_o;
  wire n3678_o;
  wire n3680_o;
  wire n3681_o;
  wire n3682_o;
  wire n3684_o;
  wire n3685_o;
  wire n3686_o;
  wire n3688_o;
  wire n3689_o;
  wire n3690_o;
  wire n3697_o;
  wire n3699_o;
  wire n3701_o;
  wire n3703_o;
  wire n3705_o;
  wire n3706_o;
  wire n3707_o;
  wire n3709_o;
  wire n3710_o;
  wire n3711_o;
  wire n3713_o;
  wire n3714_o;
  wire n3715_o;
  wire n3717_o;
  wire n3718_o;
  wire n3719_o;
  wire n3721_o;
  wire n3722_o;
  wire n3723_o;
  wire n3725_o;
  wire n3726_o;
  wire n3727_o;
  wire n3729_o;
  wire n3730_o;
  wire n3731_o;
  wire n3733_o;
  wire n3734_o;
  wire n3735_o;
  wire n3737_o;
  wire n3738_o;
  wire n3739_o;
  wire n3741_o;
  wire n3742_o;
  wire n3743_o;
  wire n3745_o;
  wire n3746_o;
  wire n3747_o;
  wire n3754_o;
  wire n3756_o;
  wire n3758_o;
  wire n3760_o;
  wire n3762_o;
  wire n3763_o;
  wire n3764_o;
  wire n3766_o;
  wire n3767_o;
  wire n3768_o;
  wire n3770_o;
  wire n3771_o;
  wire n3772_o;
  wire n3774_o;
  wire n3775_o;
  wire n3776_o;
  wire n3778_o;
  wire n3779_o;
  wire n3780_o;
  wire n3782_o;
  wire n3783_o;
  wire n3784_o;
  wire n3786_o;
  wire n3787_o;
  wire n3788_o;
  wire n3790_o;
  wire n3791_o;
  wire n3792_o;
  wire n3794_o;
  wire n3795_o;
  wire n3796_o;
  wire n3798_o;
  wire n3799_o;
  wire n3800_o;
  wire n3802_o;
  wire n3803_o;
  wire n3804_o;
  wire n3811_o;
  wire n3813_o;
  wire n3815_o;
  wire n3817_o;
  wire n3819_o;
  wire n3820_o;
  wire n3821_o;
  wire n3823_o;
  wire n3824_o;
  wire n3825_o;
  wire n3827_o;
  wire n3828_o;
  wire n3829_o;
  wire n3831_o;
  wire n3832_o;
  wire n3833_o;
  wire n3835_o;
  wire n3836_o;
  wire n3837_o;
  wire n3839_o;
  wire n3840_o;
  wire n3841_o;
  wire n3843_o;
  wire n3844_o;
  wire n3845_o;
  wire n3847_o;
  wire n3848_o;
  wire n3849_o;
  wire n3851_o;
  wire n3852_o;
  wire n3853_o;
  wire n3855_o;
  wire n3856_o;
  wire n3857_o;
  wire n3859_o;
  wire n3860_o;
  wire n3861_o;
  wire n3868_o;
  wire n3870_o;
  wire n3872_o;
  wire n3874_o;
  wire n3876_o;
  wire n3877_o;
  wire n3878_o;
  wire n3880_o;
  wire n3881_o;
  wire n3882_o;
  wire n3884_o;
  wire n3885_o;
  wire n3886_o;
  wire n3888_o;
  wire n3889_o;
  wire n3890_o;
  wire n3892_o;
  wire n3893_o;
  wire n3894_o;
  wire n3896_o;
  wire n3897_o;
  wire n3898_o;
  wire n3900_o;
  wire n3901_o;
  wire n3902_o;
  wire n3904_o;
  wire n3905_o;
  wire n3906_o;
  wire n3908_o;
  wire n3909_o;
  wire n3910_o;
  wire n3912_o;
  wire n3913_o;
  wire n3914_o;
  wire n3916_o;
  wire n3917_o;
  wire n3918_o;
  wire n3925_o;
  wire n3927_o;
  wire n3929_o;
  wire n3931_o;
  wire n3933_o;
  wire n3934_o;
  wire n3935_o;
  wire n3937_o;
  wire n3938_o;
  wire n3939_o;
  wire n3941_o;
  wire n3942_o;
  wire n3943_o;
  wire n3945_o;
  wire n3946_o;
  wire n3947_o;
  wire n3949_o;
  wire n3950_o;
  wire n3951_o;
  wire n3953_o;
  wire n3954_o;
  wire n3955_o;
  wire n3957_o;
  wire n3958_o;
  wire n3959_o;
  wire n3961_o;
  wire n3962_o;
  wire n3963_o;
  wire n3965_o;
  wire n3966_o;
  wire n3967_o;
  wire n3969_o;
  wire n3970_o;
  wire n3971_o;
  wire n3973_o;
  wire n3974_o;
  wire n3975_o;
  wire n3982_o;
  wire n3984_o;
  wire n3986_o;
  wire n3988_o;
  wire n3990_o;
  wire n3991_o;
  wire n3992_o;
  wire n3994_o;
  wire n3995_o;
  wire n3996_o;
  wire n3998_o;
  wire n3999_o;
  wire n4000_o;
  wire n4002_o;
  wire n4003_o;
  wire n4004_o;
  wire n4006_o;
  wire n4007_o;
  wire n4008_o;
  wire n4010_o;
  wire n4011_o;
  wire n4012_o;
  wire n4014_o;
  wire n4015_o;
  wire n4016_o;
  wire n4018_o;
  wire n4019_o;
  wire n4020_o;
  wire n4022_o;
  wire n4023_o;
  wire n4024_o;
  wire n4026_o;
  wire n4027_o;
  wire n4028_o;
  wire n4030_o;
  wire n4031_o;
  wire n4032_o;
  wire n4039_o;
  wire n4041_o;
  wire n4043_o;
  wire n4045_o;
  wire n4047_o;
  wire n4048_o;
  wire n4049_o;
  wire n4051_o;
  wire n4052_o;
  wire n4053_o;
  wire n4055_o;
  wire n4056_o;
  wire n4057_o;
  wire n4059_o;
  wire n4060_o;
  wire n4061_o;
  wire n4063_o;
  wire n4064_o;
  wire n4065_o;
  wire n4067_o;
  wire n4068_o;
  wire n4069_o;
  wire n4071_o;
  wire n4072_o;
  wire n4073_o;
  wire n4075_o;
  wire n4076_o;
  wire n4077_o;
  wire n4079_o;
  wire n4080_o;
  wire n4081_o;
  wire n4083_o;
  wire n4084_o;
  wire n4085_o;
  wire n4087_o;
  wire n4088_o;
  wire n4089_o;
  wire n4096_o;
  wire n4098_o;
  wire n4100_o;
  wire n4102_o;
  wire n4104_o;
  wire n4105_o;
  wire n4106_o;
  wire n4108_o;
  wire n4109_o;
  wire n4110_o;
  wire n4112_o;
  wire n4113_o;
  wire n4114_o;
  wire n4116_o;
  wire n4117_o;
  wire n4118_o;
  wire n4120_o;
  wire n4121_o;
  wire n4122_o;
  wire n4124_o;
  wire n4125_o;
  wire n4126_o;
  wire n4128_o;
  wire n4129_o;
  wire n4130_o;
  wire n4132_o;
  wire n4133_o;
  wire n4134_o;
  wire n4136_o;
  wire n4137_o;
  wire n4138_o;
  wire n4140_o;
  wire n4141_o;
  wire n4142_o;
  wire n4144_o;
  wire n4145_o;
  wire n4146_o;
  wire n4153_o;
  wire n4155_o;
  wire n4157_o;
  wire n4159_o;
  wire n4161_o;
  wire n4162_o;
  wire n4163_o;
  wire n4165_o;
  wire n4166_o;
  wire n4167_o;
  wire n4169_o;
  wire n4170_o;
  wire n4171_o;
  wire n4173_o;
  wire n4174_o;
  wire n4175_o;
  wire n4177_o;
  wire n4178_o;
  wire n4179_o;
  wire n4181_o;
  wire n4182_o;
  wire n4183_o;
  wire n4185_o;
  wire n4186_o;
  wire n4187_o;
  wire n4189_o;
  wire n4190_o;
  wire n4191_o;
  wire n4193_o;
  wire n4194_o;
  wire n4195_o;
  wire n4197_o;
  wire n4198_o;
  wire n4199_o;
  wire n4201_o;
  wire n4202_o;
  wire n4203_o;
  wire [3:0] n4204_o;
  wire [3:0] n4205_o;
  wire [3:0] n4206_o;
  wire [3:0] n4207_o;
  wire [3:0] n4208_o;
  wire [3:0] n4209_o;
  wire [3:0] n4210_o;
  wire [3:0] n4211_o;
  wire [3:0] n4212_o;
  wire [15:0] n4213_o;
  wire [15:0] n4214_o;
  wire [4:0] n4215_o;
  wire [36:0] n4216_o;
  wire n4217_o;
  wire n4218_o;
  wire n4219_o;
  wire n4220_o;
  wire n4221_o;
  wire n4222_o;
  wire n4223_o;
  wire n4224_o;
  wire n4225_o;
  wire n4226_o;
  wire n4227_o;
  wire n4228_o;
  wire n4229_o;
  wire n4230_o;
  wire n4231_o;
  wire n4232_o;
  wire n4233_o;
  wire n4234_o;
  wire n4235_o;
  wire n4236_o;
  wire n4237_o;
  wire n4238_o;
  wire n4239_o;
  wire n4240_o;
  wire n4241_o;
  wire n4242_o;
  wire n4243_o;
  wire n4244_o;
  wire n4245_o;
  wire n4246_o;
  wire n4247_o;
  wire n4248_o;
  wire n4249_o;
  wire n4250_o;
  wire n4251_o;
  wire n4252_o;
  wire n4259_o;
  wire n4261_o;
  wire n4263_o;
  wire n4265_o;
  wire n4267_o;
  wire n4268_o;
  wire n4269_o;
  wire n4271_o;
  wire n4272_o;
  wire n4273_o;
  wire n4275_o;
  wire n4276_o;
  wire n4277_o;
  wire n4279_o;
  wire n4280_o;
  wire n4281_o;
  wire n4283_o;
  wire n4284_o;
  wire n4285_o;
  wire n4287_o;
  wire n4288_o;
  wire n4289_o;
  wire n4291_o;
  wire n4292_o;
  wire n4293_o;
  wire n4295_o;
  wire n4296_o;
  wire n4297_o;
  wire n4299_o;
  wire n4300_o;
  wire n4301_o;
  wire n4303_o;
  wire n4304_o;
  wire n4305_o;
  wire n4307_o;
  wire n4308_o;
  wire n4309_o;
  wire n4311_o;
  wire n4312_o;
  wire n4313_o;
  wire n4315_o;
  wire n4316_o;
  wire n4317_o;
  wire n4319_o;
  wire n4320_o;
  wire n4321_o;
  wire n4323_o;
  wire n4324_o;
  wire n4325_o;
  wire n4327_o;
  wire n4328_o;
  wire n4329_o;
  wire n4331_o;
  wire n4332_o;
  wire n4333_o;
  wire n4335_o;
  wire n4336_o;
  wire n4337_o;
  wire n4339_o;
  wire n4340_o;
  wire n4341_o;
  wire n4343_o;
  wire n4344_o;
  wire n4345_o;
  wire n4347_o;
  wire n4348_o;
  wire n4349_o;
  wire n4351_o;
  wire n4352_o;
  wire n4353_o;
  wire n4355_o;
  wire n4356_o;
  wire n4357_o;
  wire n4359_o;
  wire n4360_o;
  wire n4361_o;
  wire n4363_o;
  wire n4364_o;
  wire n4365_o;
  wire n4367_o;
  wire n4368_o;
  wire n4369_o;
  wire n4371_o;
  wire n4372_o;
  wire n4373_o;
  wire n4375_o;
  wire n4376_o;
  wire n4377_o;
  wire n4379_o;
  wire n4380_o;
  wire n4381_o;
  wire n4383_o;
  wire n4384_o;
  wire n4385_o;
  wire n4387_o;
  wire n4388_o;
  wire n4389_o;
  wire n4391_o;
  wire n4392_o;
  wire n4393_o;
  wire n4395_o;
  wire n4396_o;
  wire n4397_o;
  wire n4399_o;
  wire n4400_o;
  wire n4401_o;
  wire n4403_o;
  wire n4404_o;
  wire n4405_o;
  wire n4412_o;
  wire n4414_o;
  wire n4416_o;
  wire n4418_o;
  wire n4420_o;
  wire n4421_o;
  wire n4422_o;
  wire n4424_o;
  wire n4425_o;
  wire n4426_o;
  wire n4428_o;
  wire n4429_o;
  wire n4430_o;
  wire n4432_o;
  wire n4433_o;
  wire n4434_o;
  wire n4436_o;
  wire n4437_o;
  wire n4438_o;
  wire n4440_o;
  wire n4441_o;
  wire n4442_o;
  wire n4444_o;
  wire n4445_o;
  wire n4446_o;
  wire n4448_o;
  wire n4449_o;
  wire n4450_o;
  wire n4452_o;
  wire n4453_o;
  wire n4454_o;
  wire n4456_o;
  wire n4457_o;
  wire n4458_o;
  wire n4460_o;
  wire n4461_o;
  wire n4462_o;
  wire n4464_o;
  wire n4465_o;
  wire n4466_o;
  wire n4468_o;
  wire n4469_o;
  wire n4470_o;
  wire n4472_o;
  wire n4473_o;
  wire n4474_o;
  wire n4476_o;
  wire n4477_o;
  wire n4478_o;
  wire n4480_o;
  wire n4481_o;
  wire n4482_o;
  wire n4484_o;
  wire n4485_o;
  wire n4486_o;
  wire n4488_o;
  wire n4489_o;
  wire n4490_o;
  wire n4492_o;
  wire n4493_o;
  wire n4494_o;
  wire n4496_o;
  wire n4497_o;
  wire n4498_o;
  wire n4500_o;
  wire n4501_o;
  wire n4502_o;
  wire n4504_o;
  wire n4505_o;
  wire n4506_o;
  wire n4508_o;
  wire n4509_o;
  wire n4510_o;
  wire n4512_o;
  wire n4513_o;
  wire n4514_o;
  wire n4516_o;
  wire n4517_o;
  wire n4518_o;
  wire n4520_o;
  wire n4521_o;
  wire n4522_o;
  wire n4524_o;
  wire n4525_o;
  wire n4526_o;
  wire n4528_o;
  wire n4529_o;
  wire n4530_o;
  wire n4532_o;
  wire n4533_o;
  wire n4534_o;
  wire n4536_o;
  wire n4537_o;
  wire n4538_o;
  wire n4540_o;
  wire n4541_o;
  wire n4542_o;
  wire n4544_o;
  wire n4545_o;
  wire n4546_o;
  wire n4548_o;
  wire n4549_o;
  wire n4550_o;
  wire n4552_o;
  wire n4553_o;
  wire n4554_o;
  wire n4556_o;
  wire n4557_o;
  wire n4558_o;
  wire n4565_o;
  wire n4567_o;
  wire n4569_o;
  wire n4571_o;
  wire n4573_o;
  wire n4574_o;
  wire n4575_o;
  wire n4577_o;
  wire n4578_o;
  wire n4579_o;
  wire n4581_o;
  wire n4582_o;
  wire n4583_o;
  wire n4585_o;
  wire n4586_o;
  wire n4587_o;
  wire n4589_o;
  wire n4590_o;
  wire n4591_o;
  wire n4593_o;
  wire n4594_o;
  wire n4595_o;
  wire n4597_o;
  wire n4598_o;
  wire n4599_o;
  wire n4601_o;
  wire n4602_o;
  wire n4603_o;
  wire n4605_o;
  wire n4606_o;
  wire n4607_o;
  wire n4609_o;
  wire n4610_o;
  wire n4611_o;
  wire n4613_o;
  wire n4614_o;
  wire n4615_o;
  wire n4617_o;
  wire n4618_o;
  wire n4619_o;
  wire n4621_o;
  wire n4622_o;
  wire n4623_o;
  wire n4625_o;
  wire n4626_o;
  wire n4627_o;
  wire n4629_o;
  wire n4630_o;
  wire n4631_o;
  wire n4633_o;
  wire n4634_o;
  wire n4635_o;
  wire n4637_o;
  wire n4638_o;
  wire n4639_o;
  wire n4641_o;
  wire n4642_o;
  wire n4643_o;
  wire n4645_o;
  wire n4646_o;
  wire n4647_o;
  wire n4649_o;
  wire n4650_o;
  wire n4651_o;
  wire n4653_o;
  wire n4654_o;
  wire n4655_o;
  wire n4657_o;
  wire n4658_o;
  wire n4659_o;
  wire n4661_o;
  wire n4662_o;
  wire n4663_o;
  wire n4665_o;
  wire n4666_o;
  wire n4667_o;
  wire n4669_o;
  wire n4670_o;
  wire n4671_o;
  wire n4673_o;
  wire n4674_o;
  wire n4675_o;
  wire n4677_o;
  wire n4678_o;
  wire n4679_o;
  wire n4681_o;
  wire n4682_o;
  wire n4683_o;
  wire n4685_o;
  wire n4686_o;
  wire n4687_o;
  wire n4689_o;
  wire n4690_o;
  wire n4691_o;
  wire n4693_o;
  wire n4694_o;
  wire n4695_o;
  wire n4697_o;
  wire n4698_o;
  wire n4699_o;
  wire n4701_o;
  wire n4702_o;
  wire n4703_o;
  wire n4705_o;
  wire n4706_o;
  wire n4707_o;
  wire n4709_o;
  wire n4710_o;
  wire n4711_o;
  wire n4718_o;
  wire n4720_o;
  wire n4722_o;
  wire n4724_o;
  wire n4726_o;
  wire n4727_o;
  wire n4728_o;
  wire n4730_o;
  wire n4731_o;
  wire n4732_o;
  wire n4734_o;
  wire n4735_o;
  wire n4736_o;
  wire n4738_o;
  wire n4739_o;
  wire n4740_o;
  wire n4742_o;
  wire n4743_o;
  wire n4744_o;
  wire n4746_o;
  wire n4747_o;
  wire n4748_o;
  wire n4750_o;
  wire n4751_o;
  wire n4752_o;
  wire n4754_o;
  wire n4755_o;
  wire n4756_o;
  wire n4758_o;
  wire n4759_o;
  wire n4760_o;
  wire n4762_o;
  wire n4763_o;
  wire n4764_o;
  wire n4766_o;
  wire n4767_o;
  wire n4768_o;
  wire n4770_o;
  wire n4771_o;
  wire n4772_o;
  wire n4774_o;
  wire n4775_o;
  wire n4776_o;
  wire n4778_o;
  wire n4779_o;
  wire n4780_o;
  wire n4782_o;
  wire n4783_o;
  wire n4784_o;
  wire n4786_o;
  wire n4787_o;
  wire n4788_o;
  wire n4790_o;
  wire n4791_o;
  wire n4792_o;
  wire n4794_o;
  wire n4795_o;
  wire n4796_o;
  wire n4798_o;
  wire n4799_o;
  wire n4800_o;
  wire n4802_o;
  wire n4803_o;
  wire n4804_o;
  wire n4806_o;
  wire n4807_o;
  wire n4808_o;
  wire n4810_o;
  wire n4811_o;
  wire n4812_o;
  wire n4814_o;
  wire n4815_o;
  wire n4816_o;
  wire n4818_o;
  wire n4819_o;
  wire n4820_o;
  wire n4822_o;
  wire n4823_o;
  wire n4824_o;
  wire n4826_o;
  wire n4827_o;
  wire n4828_o;
  wire n4830_o;
  wire n4831_o;
  wire n4832_o;
  wire n4834_o;
  wire n4835_o;
  wire n4836_o;
  wire n4838_o;
  wire n4839_o;
  wire n4840_o;
  wire n4842_o;
  wire n4843_o;
  wire n4844_o;
  wire n4846_o;
  wire n4847_o;
  wire n4848_o;
  wire n4850_o;
  wire n4851_o;
  wire n4852_o;
  wire n4854_o;
  wire n4855_o;
  wire n4856_o;
  wire n4858_o;
  wire n4859_o;
  wire n4860_o;
  wire n4862_o;
  wire n4863_o;
  wire n4864_o;
  wire n4871_o;
  wire n4873_o;
  wire n4875_o;
  wire n4877_o;
  wire n4879_o;
  wire n4880_o;
  wire n4881_o;
  wire n4883_o;
  wire n4884_o;
  wire n4885_o;
  wire n4887_o;
  wire n4888_o;
  wire n4889_o;
  wire n4891_o;
  wire n4892_o;
  wire n4893_o;
  wire n4895_o;
  wire n4896_o;
  wire n4897_o;
  wire n4899_o;
  wire n4900_o;
  wire n4901_o;
  wire n4903_o;
  wire n4904_o;
  wire n4905_o;
  wire n4907_o;
  wire n4908_o;
  wire n4909_o;
  wire n4911_o;
  wire n4912_o;
  wire n4913_o;
  wire n4915_o;
  wire n4916_o;
  wire n4917_o;
  wire n4919_o;
  wire n4920_o;
  wire n4921_o;
  wire n4923_o;
  wire n4924_o;
  wire n4925_o;
  wire n4927_o;
  wire n4928_o;
  wire n4929_o;
  wire n4931_o;
  wire n4932_o;
  wire n4933_o;
  wire n4935_o;
  wire n4936_o;
  wire n4937_o;
  wire n4939_o;
  wire n4940_o;
  wire n4941_o;
  wire n4943_o;
  wire n4944_o;
  wire n4945_o;
  wire n4947_o;
  wire n4948_o;
  wire n4949_o;
  wire n4951_o;
  wire n4952_o;
  wire n4953_o;
  wire n4955_o;
  wire n4956_o;
  wire n4957_o;
  wire n4959_o;
  wire n4960_o;
  wire n4961_o;
  wire n4963_o;
  wire n4964_o;
  wire n4965_o;
  wire n4967_o;
  wire n4968_o;
  wire n4969_o;
  wire n4971_o;
  wire n4972_o;
  wire n4973_o;
  wire n4975_o;
  wire n4976_o;
  wire n4977_o;
  wire n4979_o;
  wire n4980_o;
  wire n4981_o;
  wire n4983_o;
  wire n4984_o;
  wire n4985_o;
  wire n4987_o;
  wire n4988_o;
  wire n4989_o;
  wire n4991_o;
  wire n4992_o;
  wire n4993_o;
  wire n4995_o;
  wire n4996_o;
  wire n4997_o;
  wire n4999_o;
  wire n5000_o;
  wire n5001_o;
  wire n5003_o;
  wire n5004_o;
  wire n5005_o;
  wire n5007_o;
  wire n5008_o;
  wire n5009_o;
  wire n5011_o;
  wire n5012_o;
  wire n5013_o;
  wire n5015_o;
  wire n5016_o;
  wire n5017_o;
  wire [3:0] n5018_o;
  wire [4:0] n5019_o;
  wire [7:0] n5021_o;
  wire n5027_o;
  wire n5029_o;
  wire n5031_o;
  wire n5032_o;
  wire n5033_o;
  wire n5034_o;
  wire n5035_o;
  wire n5036_o;
  wire n5037_o;
  wire n5038_o;
  wire n5039_o;
  wire n5040_o;
  wire n5041_o;
  wire n5042_o;
  wire n5043_o;
  wire n5044_o;
  wire n5045_o;
  wire [4:0] n5046_o;
  wire [35:0] n5047_o;
  reg [4:0] cntdown_block_cntq;
  wire n5056_o;
  wire n5058_o;
  wire n5060_o;
  wire [3:0] n5061_o;
  wire n5063_o;
  wire [4:0] n5065_o;
  wire [4:0] n5066_o;
  wire [4:0] n5067_o;
  wire [4:0] n5068_o;
  wire n5073_o;
  wire n5074_o;
  wire [4:0] n5076_o;
  reg [4:0] n5077_q;
  reg [7:0] din_block_dinlat;
  wire din_block_ndincom;
  wire [7:0] din_block_latchhq;
  wire [7:0] din_block_latchh;
  wire n5081_o;
  wire n5083_o;
  wire [7:0] n5088_o;
  wire [7:0] n5089_o;
  wire n5095_o;
  wire n5097_o;
  wire n5099_o;
  wire n5100_o;
  wire n5101_o;
  wire n5102_o;
  wire n5103_o;
  wire n5104_o;
  wire n5105_o;
  wire n5106_o;
  wire n5107_o;
  wire n5108_o;
  wire n5109_o;
  wire n5110_o;
  wire n5111_o;
  wire n5112_o;
  wire n5113_o;
  wire n5121_o;
  wire n5123_o;
  wire n5125_o;
  wire [6:0] n5126_o;
  wire [7:0] n5127_o;
  wire n5134_o;
  wire n5139_o;
  wire n5140_o;
  wire n5141_o;
  wire [6:0] n5143_o;
  wire [6:0] n5144_o;
  wire n5152_o;
  wire n5154_o;
  wire n5156_o;
  wire n5157_o;
  wire n5158_o;
  wire n5159_o;
  wire [6:0] n5160_o;
  wire [15:0] n5162_o;
  wire [15:0] n5163_o;
  wire [15:0] n5164_o;
  wire [15:0] n5165_o;
  wire [7:0] n5168_o;
  reg [7:0] n5169_q;
  wire [7:0] n5170_o;
  reg [7:0] n5171_q;
  wire [7:0] n5172_o;
  reg [9:0] random_block_lfsr;
  wire random_block_all0;
  wire random_block_feedback;
  wire [8:0] n5175_o;
  wire n5181_o;
  wire n5183_o;
  wire n5185_o;
  wire n5186_o;
  wire n5187_o;
  wire n5188_o;
  wire n5189_o;
  wire n5190_o;
  wire n5191_o;
  wire n5192_o;
  wire n5193_o;
  wire n5194_o;
  wire n5195_o;
  wire n5196_o;
  wire n5197_o;
  wire n5198_o;
  wire n5199_o;
  wire n5200_o;
  wire n5201_o;
  wire n5202_o;
  wire n5203_o;
  wire n5204_o;
  wire n5205_o;
  wire n5213_o;
  wire n5215_o;
  wire [8:0] n5217_o;
  wire n5218_o;
  wire [9:0] n5219_o;
  wire n5222_o;
  wire [9:0] n5223_o;
  reg [9:0] n5224_q;
  wire start_block_nvcu;
  wire [2:0] start_block_startq;
  wire start_block_startriseq;
  wire start_block_startriseqvcu;
  wire start_block_ffsset;
  wire start_block_ffsloop;
  reg start_block_ffs1q;
  reg start_block_ffs2q;
  reg start_block_ffs3q;
  reg start_block_ffs4q;
  wire start_block_ffs1nq;
  wire start_block_ffs2nq;
  wire start_block_ffs3nq;
  wire start_block_ffs4nq;
  reg start_block_ffs5q;
  wire start_block_ffs5nq;
  wire start_block_vcumode;
  wire start_block_vcufinal;
  wire start_block_vcufinal1q;
  wire start_block_vcufinal2q;
  wire start_block_nvcufinal12;
  wire start_block_xromdo7nqdel;
  reg start_block_msff1q;
  reg start_block_msff2q;
  reg start_block_pmsff3q;
  wire start_block_msff1nq;
  wire start_block_msff2nq;
  wire start_block_pmsff3nq;
  wire start_block_msffset;
  wire start_block_n001x;
  wire start_block_n002x;
  wire start_block_n003x;
  wire start_block_n004x;
  wire start_block_n005x;
  wire start_block_n006x;
  wire start_block_n007x;
  wire start_block_n008x;
  wire start_block_n009x;
  wire start_block_n014x;
  wire start_block_n015x;
  wire start_block_n016x;
  wire start_block_n017x;
  wire [3:0] start_block_n012x;
  wire start_block_busy1q;
  wire start_block_busy2q;
  wire start_block_setbusy1;
  wire n5233_o;
  wire n5234_o;
  wire n5235_o;
  wire n5243_o;
  wire n5245_o;
  wire [1:0] n5247_o;
  wire [2:0] n5248_o;
  wire n5249_o;
  wire n5257_o;
  wire n5258_o;
  wire n5259_o;
  wire n5260_o;
  wire n5261_o;
  wire n5262_o;
  wire n5270_o;
  wire n5272_o;
  wire n5274_o;
  wire n5275_o;
  wire n5276_o;
  wire n5277_o;
  wire n5278_o;
  wire n5279_o;
  wire n5280_o;
  wire n5281_o;
  wire n5282_o;
  wire n5283_o;
  wire n5284_o;
  wire n5304_o;
  wire n5306_o;
  wire n5310_o;
  wire n5311_o;
  wire n5312_o;
  wire n5313_o;
  wire n5314_o;
  wire n5315_o;
  wire n5316_o;
  wire n5317_o;
  wire n5318_o;
  wire n5319_o;
  wire n5327_o;
  wire n5329_o;
  wire n5330_o;
  wire n5331_o;
  wire n5332_o;
  wire n5341_o;
  wire n5342_o;
  wire n5343_o;
  wire n5344_o;
  wire n5345_o;
  wire n5346_o;
  wire n5347_o;
  wire n5348_o;
  wire n5349_o;
  wire n5350_o;
  wire n5351_o;
  wire n5352_o;
  wire n5353_o;
  wire n5354_o;
  wire n5355_o;
  wire start_block_xromdo7nqdel_b_o_out;
  wire n5356_o;
  wire n5357_o;
  wire n5358_o;
  wire n5359_o;
  wire n5361_o;
  wire n5362_o;
  wire n5363_o;
  wire n5364_o;
  wire n5365_o;
  wire n5366_o;
  wire n5367_o;
  wire n5368_o;
  wire n5369_o;
  wire n5377_o;
  wire n5379_o;
  wire n5381_o;
  wire n5382_o;
  wire n5383_o;
  wire n5388_o;
  wire n5396_o;
  wire n5398_o;
  wire n5400_o;
  wire n5401_o;
  wire n5402_o;
  wire n5403_o;
  wire n5408_o;
  wire n5416_o;
  wire n5418_o;
  wire n5420_o;
  wire n5421_o;
  wire n5422_o;
  wire n5423_o;
  wire n5426_o;
  wire n5427_o;
  wire n5428_o;
  wire n5429_o;
  wire n5430_o;
  wire n5431_o;
  wire n5432_o;
  wire n5433_o;
  wire n5434_o;
  wire n5435_o;
  wire n5436_o;
  wire n5437_o;
  wire n5438_o;
  wire n5439_o;
  wire n5440_o;
  wire n5441_o;
  wire n5442_o;
  wire n5443_o;
  wire n5445_o;
  wire n5450_o;
  wire n5451_o;
  wire n5452_o;
  wire n5453_o;
  wire n5454_o;
  wire n5455_o;
  wire n5456_o;
  wire n5457_o;
  wire n5458_o;
  wire n5459_o;
  wire n5460_o;
  wire n5461_o;
  wire n5462_o;
  wire n5463_o;
  wire n5464_o;
  wire n5465_o;
  wire n5466_o;
  wire n5467_o;
  wire n5468_o;
  wire n5469_o;
  wire n5470_o;
  wire n5479_o;
  wire n5480_o;
  wire n5481_o;
  wire n5482_o;
  wire n5483_o;
  wire n5484_o;
  wire n5485_o;
  wire n5486_o;
  wire n5487_o;
  wire [3:0] n5488_o;
  wire n5493_o;
  wire n5494_o;
  wire n5495_o;
  wire n5496_o;
  wire n5497_o;
  wire n5498_o;
  wire n5499_o;
  wire n5500_o;
  wire n5501_o;
  wire [3:0] n5502_o;
  wire n5507_o;
  wire n5508_o;
  wire n5509_o;
  wire n5510_o;
  wire n5511_o;
  wire n5512_o;
  wire n5513_o;
  wire n5514_o;
  wire n5515_o;
  wire [3:0] n5516_o;
  wire n5521_o;
  wire n5522_o;
  wire n5523_o;
  wire n5524_o;
  wire n5525_o;
  wire [3:0] n5526_o;
  wire n5527_o;
  wire n5528_o;
  wire n5529_o;
  wire n5530_o;
  wire n5531_o;
  wire n5532_o;
  wire n5533_o;
  wire n5534_o;
  wire n5535_o;
  wire n5536_o;
  wire n5537_o;
  wire n5538_o;
  wire n5539_o;
  wire n5540_o;
  wire n5541_o;
  wire n5542_o;
  wire n5543_o;
  wire n5544_o;
  wire n5545_o;
  wire n5546_o;
  wire n5547_o;
  wire n5548_o;
  wire n5549_o;
  wire n5550_o;
  wire n5551_o;
  wire n5552_o;
  wire n5553_o;
  wire n5554_o;
  wire n5555_o;
  wire n5556_o;
  wire n5557_o;
  wire n5558_o;
  wire n5559_o;
  wire n5560_o;
  wire n5567_o;
  wire n5568_o;
  wire n5569_o;
  wire n5570_o;
  wire n5571_o;
  wire n5572_o;
  wire n5573_o;
  wire [3:0] n5574_o;
  wire n5576_o;
  wire n5577_o;
  wire n5582_o;
  wire n5583_o;
  wire n5584_o;
  wire n5585_o;
  wire n5586_o;
  wire n5587_o;
  wire n5588_o;
  wire [3:0] n5589_o;
  wire n5594_o;
  wire n5595_o;
  wire n5596_o;
  wire n5597_o;
  wire n5598_o;
  wire n5599_o;
  wire n5600_o;
  wire n5601_o;
  wire n5602_o;
  wire n5603_o;
  wire n5604_o;
  wire n5605_o;
  wire n5606_o;
  wire n5607_o;
  wire n5608_o;
  wire n5609_o;
  wire n5610_o;
  wire n5611_o;
  wire n5612_o;
  wire n5613_o;
  wire n5614_o;
  wire n5615_o;
  wire n5616_o;
  wire n5617_o;
  wire n5618_o;
  wire n5619_o;
  wire n5620_o;
  wire n5621_o;
  wire [3:0] n5622_o;
  wire n5628_o;
  wire n5629_o;
  wire n5630_o;
  wire n5631_o;
  wire n5632_o;
  wire n5640_o;
  wire n5642_o;
  wire n5644_o;
  wire n5645_o;
  wire n5657_o;
  wire n5659_o;
  wire n5661_o;
  wire n5662_o;
  wire n5667_o;
  wire n5668_o;
  wire n5669_o;
  wire n5670_o;
  wire n5671_o;
  wire n5672_o;
  wire n5674_o;
  wire n5679_o;
  wire n5680_o;
  wire n5681_o;
  wire n5682_o;
  wire n5683_o;
  wire n5684_o;
  wire n5685_o;
  wire n5686_o;
  wire n5687_o;
  wire n5688_o;
  wire n5689_o;
  wire n5690_o;
  wire n5691_o;
  wire n5692_o;
  wire n5693_o;
  wire n5695_o;
  wire n5696_o;
  wire n5697_o;
  wire n5702_o;
  wire n5703_o;
  wire n5704_o;
  wire n5711_o;
  wire n5712_o;
  wire n5717_o;
  wire n5718_o;
  wire n5719_o;
  wire n5720_o;
  wire [2:0] n5721_o;
  reg [2:0] n5722_q;
  wire n5723_o;
  reg n5724_q;
  wire n5725_o;
  reg n5726_q;
  wire n5727_o;
  wire n5728_o;
  wire n5729_o;
  reg n5730_q;
  wire n5731_o;
  reg n5732_q;
  wire n5733_o;
  reg n5734_q;
  wire n5735_o;
  reg n5736_q;
  wire n5737_o;
  reg n5738_q;
  wire n5739_o;
  reg n5740_q;
  wire n5741_o;
  reg n5742_q;
  wire n5743_o;
  reg n5744_q;
  wire n5745_o;
  reg n5746_q;
  wire n5747_o;
  reg n5748_q;
  wire n5749_o;
  reg n5750_q;
  wire [4:0] krom_block_ka;
  wire krom_block_agen_block_nfsrdo6;
  wire [3:0] krom_block_agen_block_ksaq;
  wire [4:0] n5751_o;
  reg [4:0] krom_block_agen_block_n5752_toggle;
  wire n5755_o;
  wire n5761_o;
  wire n5763_o;
  wire [3:0] n5766_o;
  wire [4:0] n5767_o;
  wire n5768_o;
  wire n5769_o;
  wire n5770_o;
  wire n5771_o;
  wire n5772_o;
  wire n5773_o;
  wire [3:0] n5774_o;
  wire [4:0] n5775_o;
  wire n5776_o;
  wire n5777_o;
  wire n5778_o;
  wire [2:0] n5779_o;
  wire [4:0] n5780_o;
  wire n5781_o;
  wire n5782_o;
  wire n5783_o;
  wire n5784_o;
  wire n5785_o;
  wire n5786_o;
  wire [2:0] n5787_o;
  wire [4:0] n5788_o;
  wire n5789_o;
  wire n5790_o;
  wire n5791_o;
  wire [1:0] n5792_o;
  wire [4:0] n5793_o;
  wire n5794_o;
  wire n5795_o;
  wire n5796_o;
  wire n5797_o;
  wire n5798_o;
  wire n5799_o;
  wire [1:0] n5800_o;
  wire [4:0] n5801_o;
  wire n5802_o;
  wire n5803_o;
  wire n5804_o;
  wire n5805_o;
  wire [4:0] n5806_o;
  wire n5807_o;
  wire n5808_o;
  wire n5809_o;
  wire n5810_o;
  wire n5811_o;
  wire n5812_o;
  wire n5813_o;
  wire [4:0] n5814_o;
  wire n5815_o;
  wire n5816_o;
  wire n5817_o;
  wire [3:0] n5818_o;
  wire [4:0] n5820_o;
  wire n5826_o;
  wire n5827_o;
  wire [4:0] n5828_o;
  reg [4:0] n5829_q;
  wire n5830_o;
  wire n5831_o;
  wire n5832_o;
  wire n5833_o;
  wire n5834_o;
  wire n5835_o;
  wire n5836_o;
  wire n5837_o;
  wire n5838_o;
  wire n5839_o;
  wire n5840_o;
  wire n5841_o;
  wire n5842_o;
  wire n5843_o;
  wire n5844_o;
  wire n5845_o;
  wire n5846_o;
  wire n5847_o;
  wire n5848_o;
  wire n5849_o;
  wire n5850_o;
  wire n5851_o;
  wire n5852_o;
  wire n5853_o;
  wire n5854_o;
  wire n5855_o;
  wire n5856_o;
  wire n5857_o;
  wire n5858_o;
  wire n5859_o;
  wire n5860_o;
  wire [3:0] n5861_o;
  wire [3:0] n5862_o;
  reg [3:0] n5863_q;
  wire [9:0] krom_block_rom_block_kslice0;
  wire [9:0] krom_block_rom_block_kslice1;
  wire [9:0] krom_block_rom_block_kslice2;
  wire [9:0] krom_block_rom_block_kslice3;
  wire [9:0] krom_block_rom_block_kslice4;
  wire [9:0] krom_block_rom_block_kslice5;
  wire [31:0] krom_block_rom_block_wl;
  wire [5:0] krom_block_rom_block_wl_slice;
  wire krom_block_rom_block_nkaodd;
  wire krom_block_rom_block_nksa0;
  wire krom_block_rom_block_range_s0s1s2;
  wire krom_block_rom_block_range_s3s4;
  wire [9:0] krom_block_rom_block_kout;
  wire [4:0] n5868_o;
  localparam [31:0] n5870_o = 32'b00000000000000000000000000000000;
  wire n5886_o;
  wire n5888_o;
  wire n5890_o;
  wire n5892_o;
  wire n5894_o;
  wire n5895_o;
  wire n5896_o;
  wire n5898_o;
  wire n5899_o;
  wire n5900_o;
  wire n5902_o;
  wire n5903_o;
  wire n5904_o;
  wire n5906_o;
  wire n5907_o;
  wire n5908_o;
  wire n5910_o;
  wire n5911_o;
  wire n5912_o;
  wire n5914_o;
  wire n5915_o;
  wire n5916_o;
  wire n5918_o;
  wire n5919_o;
  wire n5920_o;
  wire n5922_o;
  wire n5923_o;
  wire n5924_o;
  wire n5926_o;
  wire n5927_o;
  wire n5928_o;
  wire n5930_o;
  wire n5931_o;
  wire n5932_o;
  wire n5934_o;
  wire n5935_o;
  wire n5936_o;
  wire n5938_o;
  wire n5939_o;
  wire n5940_o;
  wire n5942_o;
  wire n5943_o;
  wire n5944_o;
  wire n5946_o;
  wire n5947_o;
  wire n5948_o;
  wire n5950_o;
  wire n5951_o;
  wire n5952_o;
  wire n5954_o;
  wire n5955_o;
  wire n5956_o;
  wire n5958_o;
  wire n5959_o;
  wire n5960_o;
  wire n5962_o;
  wire n5963_o;
  wire n5964_o;
  wire n5966_o;
  wire n5967_o;
  wire n5968_o;
  wire n5970_o;
  wire n5971_o;
  wire n5972_o;
  wire n5974_o;
  wire n5975_o;
  wire n5976_o;
  wire n5978_o;
  wire n5979_o;
  wire n5980_o;
  wire n5982_o;
  wire n5983_o;
  wire n5984_o;
  wire n5986_o;
  wire n5987_o;
  wire n5988_o;
  wire n5990_o;
  wire n5991_o;
  wire n5992_o;
  wire n5994_o;
  wire n5995_o;
  wire n5996_o;
  wire n5998_o;
  wire n5999_o;
  wire n6000_o;
  wire n6002_o;
  wire n6003_o;
  wire n6004_o;
  wire n6006_o;
  wire n6007_o;
  wire n6008_o;
  wire n6010_o;
  wire n6011_o;
  wire n6012_o;
  wire n6014_o;
  wire n6015_o;
  wire n6016_o;
  wire n6017_o;
  wire n6029_o;
  wire n6031_o;
  wire n6033_o;
  wire n6035_o;
  wire n6037_o;
  wire n6038_o;
  wire n6039_o;
  wire n6041_o;
  wire n6042_o;
  wire n6043_o;
  wire n6045_o;
  wire n6046_o;
  wire n6047_o;
  wire n6049_o;
  wire n6050_o;
  wire n6051_o;
  wire n6053_o;
  wire n6054_o;
  wire n6055_o;
  wire n6057_o;
  wire n6058_o;
  wire n6059_o;
  wire n6061_o;
  wire n6062_o;
  wire n6063_o;
  wire n6065_o;
  wire n6066_o;
  wire n6067_o;
  wire n6069_o;
  wire n6070_o;
  wire n6071_o;
  wire n6073_o;
  wire n6074_o;
  wire n6075_o;
  wire n6077_o;
  wire n6078_o;
  wire n6079_o;
  wire n6081_o;
  wire n6082_o;
  wire n6083_o;
  wire n6085_o;
  wire n6086_o;
  wire n6087_o;
  wire n6089_o;
  wire n6090_o;
  wire n6091_o;
  wire n6093_o;
  wire n6094_o;
  wire n6095_o;
  wire n6097_o;
  wire n6098_o;
  wire n6099_o;
  wire n6101_o;
  wire n6102_o;
  wire n6103_o;
  wire n6105_o;
  wire n6106_o;
  wire n6107_o;
  wire n6109_o;
  wire n6110_o;
  wire n6111_o;
  wire n6113_o;
  wire n6114_o;
  wire n6115_o;
  wire n6117_o;
  wire n6118_o;
  wire n6119_o;
  wire n6121_o;
  wire n6122_o;
  wire n6123_o;
  wire n6125_o;
  wire n6126_o;
  wire n6127_o;
  wire n6129_o;
  wire n6130_o;
  wire n6131_o;
  wire n6133_o;
  wire n6134_o;
  wire n6135_o;
  wire n6137_o;
  wire n6138_o;
  wire n6139_o;
  wire n6141_o;
  wire n6142_o;
  wire n6143_o;
  wire n6145_o;
  wire n6146_o;
  wire n6147_o;
  wire n6149_o;
  wire n6150_o;
  wire n6151_o;
  wire n6153_o;
  wire n6154_o;
  wire n6155_o;
  wire n6157_o;
  wire n6158_o;
  wire n6159_o;
  wire n6160_o;
  wire n6172_o;
  wire n6174_o;
  wire n6176_o;
  wire n6178_o;
  wire n6180_o;
  wire n6181_o;
  wire n6182_o;
  wire n6184_o;
  wire n6185_o;
  wire n6186_o;
  wire n6188_o;
  wire n6189_o;
  wire n6190_o;
  wire n6192_o;
  wire n6193_o;
  wire n6194_o;
  wire n6196_o;
  wire n6197_o;
  wire n6198_o;
  wire n6200_o;
  wire n6201_o;
  wire n6202_o;
  wire n6204_o;
  wire n6205_o;
  wire n6206_o;
  wire n6208_o;
  wire n6209_o;
  wire n6210_o;
  wire n6212_o;
  wire n6213_o;
  wire n6214_o;
  wire n6216_o;
  wire n6217_o;
  wire n6218_o;
  wire n6220_o;
  wire n6221_o;
  wire n6222_o;
  wire n6224_o;
  wire n6225_o;
  wire n6226_o;
  wire n6228_o;
  wire n6229_o;
  wire n6230_o;
  wire n6232_o;
  wire n6233_o;
  wire n6234_o;
  wire n6236_o;
  wire n6237_o;
  wire n6238_o;
  wire n6240_o;
  wire n6241_o;
  wire n6242_o;
  wire n6244_o;
  wire n6245_o;
  wire n6246_o;
  wire n6248_o;
  wire n6249_o;
  wire n6250_o;
  wire n6252_o;
  wire n6253_o;
  wire n6254_o;
  wire n6256_o;
  wire n6257_o;
  wire n6258_o;
  wire n6260_o;
  wire n6261_o;
  wire n6262_o;
  wire n6264_o;
  wire n6265_o;
  wire n6266_o;
  wire n6268_o;
  wire n6269_o;
  wire n6270_o;
  wire n6272_o;
  wire n6273_o;
  wire n6274_o;
  wire n6276_o;
  wire n6277_o;
  wire n6278_o;
  wire n6280_o;
  wire n6281_o;
  wire n6282_o;
  wire n6284_o;
  wire n6285_o;
  wire n6286_o;
  wire n6288_o;
  wire n6289_o;
  wire n6290_o;
  wire n6292_o;
  wire n6293_o;
  wire n6294_o;
  wire n6296_o;
  wire n6297_o;
  wire n6298_o;
  wire n6300_o;
  wire n6301_o;
  wire n6302_o;
  wire n6303_o;
  wire n6315_o;
  wire n6317_o;
  wire n6319_o;
  wire n6321_o;
  wire n6323_o;
  wire n6324_o;
  wire n6325_o;
  wire n6327_o;
  wire n6328_o;
  wire n6329_o;
  wire n6331_o;
  wire n6332_o;
  wire n6333_o;
  wire n6335_o;
  wire n6336_o;
  wire n6337_o;
  wire n6339_o;
  wire n6340_o;
  wire n6341_o;
  wire n6343_o;
  wire n6344_o;
  wire n6345_o;
  wire n6347_o;
  wire n6348_o;
  wire n6349_o;
  wire n6351_o;
  wire n6352_o;
  wire n6353_o;
  wire n6355_o;
  wire n6356_o;
  wire n6357_o;
  wire n6359_o;
  wire n6360_o;
  wire n6361_o;
  wire n6363_o;
  wire n6364_o;
  wire n6365_o;
  wire n6367_o;
  wire n6368_o;
  wire n6369_o;
  wire n6371_o;
  wire n6372_o;
  wire n6373_o;
  wire n6375_o;
  wire n6376_o;
  wire n6377_o;
  wire n6379_o;
  wire n6380_o;
  wire n6381_o;
  wire n6383_o;
  wire n6384_o;
  wire n6385_o;
  wire n6387_o;
  wire n6388_o;
  wire n6389_o;
  wire n6391_o;
  wire n6392_o;
  wire n6393_o;
  wire n6395_o;
  wire n6396_o;
  wire n6397_o;
  wire n6399_o;
  wire n6400_o;
  wire n6401_o;
  wire n6403_o;
  wire n6404_o;
  wire n6405_o;
  wire n6407_o;
  wire n6408_o;
  wire n6409_o;
  wire n6411_o;
  wire n6412_o;
  wire n6413_o;
  wire n6415_o;
  wire n6416_o;
  wire n6417_o;
  wire n6419_o;
  wire n6420_o;
  wire n6421_o;
  wire n6423_o;
  wire n6424_o;
  wire n6425_o;
  wire n6427_o;
  wire n6428_o;
  wire n6429_o;
  wire n6431_o;
  wire n6432_o;
  wire n6433_o;
  wire n6435_o;
  wire n6436_o;
  wire n6437_o;
  wire n6439_o;
  wire n6440_o;
  wire n6441_o;
  wire n6443_o;
  wire n6444_o;
  wire n6445_o;
  wire n6446_o;
  wire n6458_o;
  wire n6460_o;
  wire n6462_o;
  wire n6464_o;
  wire n6466_o;
  wire n6467_o;
  wire n6468_o;
  wire n6470_o;
  wire n6471_o;
  wire n6472_o;
  wire n6474_o;
  wire n6475_o;
  wire n6476_o;
  wire n6478_o;
  wire n6479_o;
  wire n6480_o;
  wire n6482_o;
  wire n6483_o;
  wire n6484_o;
  wire n6486_o;
  wire n6487_o;
  wire n6488_o;
  wire n6490_o;
  wire n6491_o;
  wire n6492_o;
  wire n6494_o;
  wire n6495_o;
  wire n6496_o;
  wire n6498_o;
  wire n6499_o;
  wire n6500_o;
  wire n6502_o;
  wire n6503_o;
  wire n6504_o;
  wire n6506_o;
  wire n6507_o;
  wire n6508_o;
  wire n6510_o;
  wire n6511_o;
  wire n6512_o;
  wire n6514_o;
  wire n6515_o;
  wire n6516_o;
  wire n6518_o;
  wire n6519_o;
  wire n6520_o;
  wire n6522_o;
  wire n6523_o;
  wire n6524_o;
  wire n6526_o;
  wire n6527_o;
  wire n6528_o;
  wire n6530_o;
  wire n6531_o;
  wire n6532_o;
  wire n6534_o;
  wire n6535_o;
  wire n6536_o;
  wire n6538_o;
  wire n6539_o;
  wire n6540_o;
  wire n6542_o;
  wire n6543_o;
  wire n6544_o;
  wire n6546_o;
  wire n6547_o;
  wire n6548_o;
  wire n6550_o;
  wire n6551_o;
  wire n6552_o;
  wire n6554_o;
  wire n6555_o;
  wire n6556_o;
  wire n6558_o;
  wire n6559_o;
  wire n6560_o;
  wire n6562_o;
  wire n6563_o;
  wire n6564_o;
  wire n6566_o;
  wire n6567_o;
  wire n6568_o;
  wire n6570_o;
  wire n6571_o;
  wire n6572_o;
  wire n6574_o;
  wire n6575_o;
  wire n6576_o;
  wire n6578_o;
  wire n6579_o;
  wire n6580_o;
  wire n6582_o;
  wire n6583_o;
  wire n6584_o;
  wire n6586_o;
  wire n6587_o;
  wire n6588_o;
  wire n6589_o;
  wire n6601_o;
  wire n6603_o;
  wire n6605_o;
  wire n6607_o;
  wire n6609_o;
  wire n6610_o;
  wire n6611_o;
  wire n6613_o;
  wire n6614_o;
  wire n6615_o;
  wire n6617_o;
  wire n6618_o;
  wire n6619_o;
  wire n6621_o;
  wire n6622_o;
  wire n6623_o;
  wire n6625_o;
  wire n6626_o;
  wire n6627_o;
  wire n6629_o;
  wire n6630_o;
  wire n6631_o;
  wire n6633_o;
  wire n6634_o;
  wire n6635_o;
  wire n6637_o;
  wire n6638_o;
  wire n6639_o;
  wire n6641_o;
  wire n6642_o;
  wire n6643_o;
  wire n6645_o;
  wire n6646_o;
  wire n6647_o;
  wire n6649_o;
  wire n6650_o;
  wire n6651_o;
  wire n6653_o;
  wire n6654_o;
  wire n6655_o;
  wire n6657_o;
  wire n6658_o;
  wire n6659_o;
  wire n6661_o;
  wire n6662_o;
  wire n6663_o;
  wire n6665_o;
  wire n6666_o;
  wire n6667_o;
  wire n6669_o;
  wire n6670_o;
  wire n6671_o;
  wire n6673_o;
  wire n6674_o;
  wire n6675_o;
  wire n6677_o;
  wire n6678_o;
  wire n6679_o;
  wire n6681_o;
  wire n6682_o;
  wire n6683_o;
  wire n6685_o;
  wire n6686_o;
  wire n6687_o;
  wire n6689_o;
  wire n6690_o;
  wire n6691_o;
  wire n6693_o;
  wire n6694_o;
  wire n6695_o;
  wire n6697_o;
  wire n6698_o;
  wire n6699_o;
  wire n6701_o;
  wire n6702_o;
  wire n6703_o;
  wire n6705_o;
  wire n6706_o;
  wire n6707_o;
  wire n6709_o;
  wire n6710_o;
  wire n6711_o;
  wire n6713_o;
  wire n6714_o;
  wire n6715_o;
  wire n6717_o;
  wire n6718_o;
  wire n6719_o;
  wire n6721_o;
  wire n6722_o;
  wire n6723_o;
  wire n6725_o;
  wire n6726_o;
  wire n6727_o;
  wire n6729_o;
  wire n6730_o;
  wire n6731_o;
  wire n6732_o;
  wire n6744_o;
  wire n6746_o;
  wire n6748_o;
  wire n6750_o;
  wire n6752_o;
  wire n6753_o;
  wire n6754_o;
  wire n6756_o;
  wire n6757_o;
  wire n6758_o;
  wire n6760_o;
  wire n6761_o;
  wire n6762_o;
  wire n6764_o;
  wire n6765_o;
  wire n6766_o;
  wire n6768_o;
  wire n6769_o;
  wire n6770_o;
  wire n6772_o;
  wire n6773_o;
  wire n6774_o;
  wire n6776_o;
  wire n6777_o;
  wire n6778_o;
  wire n6780_o;
  wire n6781_o;
  wire n6782_o;
  wire n6784_o;
  wire n6785_o;
  wire n6786_o;
  wire n6788_o;
  wire n6789_o;
  wire n6790_o;
  wire n6792_o;
  wire n6793_o;
  wire n6794_o;
  wire n6796_o;
  wire n6797_o;
  wire n6798_o;
  wire n6800_o;
  wire n6801_o;
  wire n6802_o;
  wire n6804_o;
  wire n6805_o;
  wire n6806_o;
  wire n6808_o;
  wire n6809_o;
  wire n6810_o;
  wire n6812_o;
  wire n6813_o;
  wire n6814_o;
  wire n6816_o;
  wire n6817_o;
  wire n6818_o;
  wire n6820_o;
  wire n6821_o;
  wire n6822_o;
  wire n6824_o;
  wire n6825_o;
  wire n6826_o;
  wire n6828_o;
  wire n6829_o;
  wire n6830_o;
  wire n6832_o;
  wire n6833_o;
  wire n6834_o;
  wire n6836_o;
  wire n6837_o;
  wire n6838_o;
  wire n6840_o;
  wire n6841_o;
  wire n6842_o;
  wire n6844_o;
  wire n6845_o;
  wire n6846_o;
  wire n6848_o;
  wire n6849_o;
  wire n6850_o;
  wire n6852_o;
  wire n6853_o;
  wire n6854_o;
  wire n6856_o;
  wire n6857_o;
  wire n6858_o;
  wire n6860_o;
  wire n6861_o;
  wire n6862_o;
  wire n6864_o;
  wire n6865_o;
  wire n6866_o;
  wire n6868_o;
  wire n6869_o;
  wire n6870_o;
  wire n6872_o;
  wire n6873_o;
  wire n6874_o;
  wire n6875_o;
  wire n6887_o;
  wire n6889_o;
  wire n6891_o;
  wire n6893_o;
  wire n6895_o;
  wire n6896_o;
  wire n6897_o;
  wire n6899_o;
  wire n6900_o;
  wire n6901_o;
  wire n6903_o;
  wire n6904_o;
  wire n6905_o;
  wire n6907_o;
  wire n6908_o;
  wire n6909_o;
  wire n6911_o;
  wire n6912_o;
  wire n6913_o;
  wire n6915_o;
  wire n6916_o;
  wire n6917_o;
  wire n6919_o;
  wire n6920_o;
  wire n6921_o;
  wire n6923_o;
  wire n6924_o;
  wire n6925_o;
  wire n6927_o;
  wire n6928_o;
  wire n6929_o;
  wire n6931_o;
  wire n6932_o;
  wire n6933_o;
  wire n6935_o;
  wire n6936_o;
  wire n6937_o;
  wire n6939_o;
  wire n6940_o;
  wire n6941_o;
  wire n6943_o;
  wire n6944_o;
  wire n6945_o;
  wire n6947_o;
  wire n6948_o;
  wire n6949_o;
  wire n6951_o;
  wire n6952_o;
  wire n6953_o;
  wire n6955_o;
  wire n6956_o;
  wire n6957_o;
  wire n6959_o;
  wire n6960_o;
  wire n6961_o;
  wire n6963_o;
  wire n6964_o;
  wire n6965_o;
  wire n6967_o;
  wire n6968_o;
  wire n6969_o;
  wire n6971_o;
  wire n6972_o;
  wire n6973_o;
  wire n6975_o;
  wire n6976_o;
  wire n6977_o;
  wire n6979_o;
  wire n6980_o;
  wire n6981_o;
  wire n6983_o;
  wire n6984_o;
  wire n6985_o;
  wire n6987_o;
  wire n6988_o;
  wire n6989_o;
  wire n6991_o;
  wire n6992_o;
  wire n6993_o;
  wire n6995_o;
  wire n6996_o;
  wire n6997_o;
  wire n6999_o;
  wire n7000_o;
  wire n7001_o;
  wire n7003_o;
  wire n7004_o;
  wire n7005_o;
  wire n7007_o;
  wire n7008_o;
  wire n7009_o;
  wire n7011_o;
  wire n7012_o;
  wire n7013_o;
  wire n7015_o;
  wire n7016_o;
  wire n7017_o;
  wire n7018_o;
  wire n7030_o;
  wire n7032_o;
  wire n7034_o;
  wire n7036_o;
  wire n7038_o;
  wire n7039_o;
  wire n7040_o;
  wire n7042_o;
  wire n7043_o;
  wire n7044_o;
  wire n7046_o;
  wire n7047_o;
  wire n7048_o;
  wire n7050_o;
  wire n7051_o;
  wire n7052_o;
  wire n7054_o;
  wire n7055_o;
  wire n7056_o;
  wire n7058_o;
  wire n7059_o;
  wire n7060_o;
  wire n7062_o;
  wire n7063_o;
  wire n7064_o;
  wire n7066_o;
  wire n7067_o;
  wire n7068_o;
  wire n7070_o;
  wire n7071_o;
  wire n7072_o;
  wire n7074_o;
  wire n7075_o;
  wire n7076_o;
  wire n7078_o;
  wire n7079_o;
  wire n7080_o;
  wire n7082_o;
  wire n7083_o;
  wire n7084_o;
  wire n7086_o;
  wire n7087_o;
  wire n7088_o;
  wire n7090_o;
  wire n7091_o;
  wire n7092_o;
  wire n7094_o;
  wire n7095_o;
  wire n7096_o;
  wire n7098_o;
  wire n7099_o;
  wire n7100_o;
  wire n7102_o;
  wire n7103_o;
  wire n7104_o;
  wire n7106_o;
  wire n7107_o;
  wire n7108_o;
  wire n7110_o;
  wire n7111_o;
  wire n7112_o;
  wire n7114_o;
  wire n7115_o;
  wire n7116_o;
  wire n7118_o;
  wire n7119_o;
  wire n7120_o;
  wire n7122_o;
  wire n7123_o;
  wire n7124_o;
  wire n7126_o;
  wire n7127_o;
  wire n7128_o;
  wire n7130_o;
  wire n7131_o;
  wire n7132_o;
  wire n7134_o;
  wire n7135_o;
  wire n7136_o;
  wire n7138_o;
  wire n7139_o;
  wire n7140_o;
  wire n7142_o;
  wire n7143_o;
  wire n7144_o;
  wire n7146_o;
  wire n7147_o;
  wire n7148_o;
  wire n7150_o;
  wire n7151_o;
  wire n7152_o;
  wire n7154_o;
  wire n7155_o;
  wire n7156_o;
  wire n7158_o;
  wire n7159_o;
  wire n7160_o;
  wire n7161_o;
  wire n7173_o;
  wire n7175_o;
  wire n7177_o;
  wire n7179_o;
  wire n7181_o;
  wire n7182_o;
  wire n7183_o;
  wire n7185_o;
  wire n7186_o;
  wire n7187_o;
  wire n7189_o;
  wire n7190_o;
  wire n7191_o;
  wire n7193_o;
  wire n7194_o;
  wire n7195_o;
  wire n7197_o;
  wire n7198_o;
  wire n7199_o;
  wire n7201_o;
  wire n7202_o;
  wire n7203_o;
  wire n7205_o;
  wire n7206_o;
  wire n7207_o;
  wire n7209_o;
  wire n7210_o;
  wire n7211_o;
  wire n7213_o;
  wire n7214_o;
  wire n7215_o;
  wire n7217_o;
  wire n7218_o;
  wire n7219_o;
  wire n7221_o;
  wire n7222_o;
  wire n7223_o;
  wire n7225_o;
  wire n7226_o;
  wire n7227_o;
  wire n7229_o;
  wire n7230_o;
  wire n7231_o;
  wire n7233_o;
  wire n7234_o;
  wire n7235_o;
  wire n7237_o;
  wire n7238_o;
  wire n7239_o;
  wire n7241_o;
  wire n7242_o;
  wire n7243_o;
  wire n7245_o;
  wire n7246_o;
  wire n7247_o;
  wire n7249_o;
  wire n7250_o;
  wire n7251_o;
  wire n7253_o;
  wire n7254_o;
  wire n7255_o;
  wire n7257_o;
  wire n7258_o;
  wire n7259_o;
  wire n7261_o;
  wire n7262_o;
  wire n7263_o;
  wire n7265_o;
  wire n7266_o;
  wire n7267_o;
  wire n7269_o;
  wire n7270_o;
  wire n7271_o;
  wire n7273_o;
  wire n7274_o;
  wire n7275_o;
  wire n7277_o;
  wire n7278_o;
  wire n7279_o;
  wire n7281_o;
  wire n7282_o;
  wire n7283_o;
  wire n7285_o;
  wire n7286_o;
  wire n7287_o;
  wire n7289_o;
  wire n7290_o;
  wire n7291_o;
  wire n7293_o;
  wire n7294_o;
  wire n7295_o;
  wire n7297_o;
  wire n7298_o;
  wire n7299_o;
  wire n7301_o;
  wire n7302_o;
  wire n7303_o;
  wire n7304_o;
  wire [3:0] n7305_o;
  wire [3:0] n7306_o;
  wire [1:0] n7307_o;
  wire [9:0] n7308_o;
  wire n7320_o;
  wire n7322_o;
  wire n7324_o;
  wire n7326_o;
  wire n7328_o;
  wire n7329_o;
  wire n7330_o;
  wire n7332_o;
  wire n7333_o;
  wire n7334_o;
  wire n7336_o;
  wire n7337_o;
  wire n7338_o;
  wire n7340_o;
  wire n7341_o;
  wire n7342_o;
  wire n7344_o;
  wire n7345_o;
  wire n7346_o;
  wire n7348_o;
  wire n7349_o;
  wire n7350_o;
  wire n7352_o;
  wire n7353_o;
  wire n7354_o;
  wire n7356_o;
  wire n7357_o;
  wire n7358_o;
  wire n7360_o;
  wire n7361_o;
  wire n7362_o;
  wire n7364_o;
  wire n7365_o;
  wire n7366_o;
  wire n7368_o;
  wire n7369_o;
  wire n7370_o;
  wire n7372_o;
  wire n7373_o;
  wire n7374_o;
  wire n7376_o;
  wire n7377_o;
  wire n7378_o;
  wire n7380_o;
  wire n7381_o;
  wire n7382_o;
  wire n7384_o;
  wire n7385_o;
  wire n7386_o;
  wire n7388_o;
  wire n7389_o;
  wire n7390_o;
  wire n7392_o;
  wire n7393_o;
  wire n7394_o;
  wire n7396_o;
  wire n7397_o;
  wire n7398_o;
  wire n7400_o;
  wire n7401_o;
  wire n7402_o;
  wire n7404_o;
  wire n7405_o;
  wire n7406_o;
  wire n7408_o;
  wire n7409_o;
  wire n7410_o;
  wire n7412_o;
  wire n7413_o;
  wire n7414_o;
  wire n7416_o;
  wire n7417_o;
  wire n7418_o;
  wire n7420_o;
  wire n7421_o;
  wire n7422_o;
  wire n7424_o;
  wire n7425_o;
  wire n7426_o;
  wire n7428_o;
  wire n7429_o;
  wire n7430_o;
  wire n7432_o;
  wire n7433_o;
  wire n7434_o;
  wire n7436_o;
  wire n7437_o;
  wire n7438_o;
  wire n7440_o;
  wire n7441_o;
  wire n7442_o;
  wire n7444_o;
  wire n7445_o;
  wire n7446_o;
  wire n7448_o;
  wire n7449_o;
  wire n7450_o;
  wire n7451_o;
  wire n7463_o;
  wire n7465_o;
  wire n7467_o;
  wire n7469_o;
  wire n7471_o;
  wire n7472_o;
  wire n7473_o;
  wire n7475_o;
  wire n7476_o;
  wire n7477_o;
  wire n7479_o;
  wire n7480_o;
  wire n7481_o;
  wire n7483_o;
  wire n7484_o;
  wire n7485_o;
  wire n7487_o;
  wire n7488_o;
  wire n7489_o;
  wire n7491_o;
  wire n7492_o;
  wire n7493_o;
  wire n7495_o;
  wire n7496_o;
  wire n7497_o;
  wire n7499_o;
  wire n7500_o;
  wire n7501_o;
  wire n7503_o;
  wire n7504_o;
  wire n7505_o;
  wire n7507_o;
  wire n7508_o;
  wire n7509_o;
  wire n7511_o;
  wire n7512_o;
  wire n7513_o;
  wire n7515_o;
  wire n7516_o;
  wire n7517_o;
  wire n7519_o;
  wire n7520_o;
  wire n7521_o;
  wire n7523_o;
  wire n7524_o;
  wire n7525_o;
  wire n7527_o;
  wire n7528_o;
  wire n7529_o;
  wire n7531_o;
  wire n7532_o;
  wire n7533_o;
  wire n7535_o;
  wire n7536_o;
  wire n7537_o;
  wire n7539_o;
  wire n7540_o;
  wire n7541_o;
  wire n7543_o;
  wire n7544_o;
  wire n7545_o;
  wire n7547_o;
  wire n7548_o;
  wire n7549_o;
  wire n7551_o;
  wire n7552_o;
  wire n7553_o;
  wire n7555_o;
  wire n7556_o;
  wire n7557_o;
  wire n7559_o;
  wire n7560_o;
  wire n7561_o;
  wire n7563_o;
  wire n7564_o;
  wire n7565_o;
  wire n7567_o;
  wire n7568_o;
  wire n7569_o;
  wire n7571_o;
  wire n7572_o;
  wire n7573_o;
  wire n7575_o;
  wire n7576_o;
  wire n7577_o;
  wire n7579_o;
  wire n7580_o;
  wire n7581_o;
  wire n7583_o;
  wire n7584_o;
  wire n7585_o;
  wire n7587_o;
  wire n7588_o;
  wire n7589_o;
  wire n7591_o;
  wire n7592_o;
  wire n7593_o;
  wire n7594_o;
  wire n7606_o;
  wire n7608_o;
  wire n7610_o;
  wire n7612_o;
  wire n7614_o;
  wire n7615_o;
  wire n7616_o;
  wire n7618_o;
  wire n7619_o;
  wire n7620_o;
  wire n7622_o;
  wire n7623_o;
  wire n7624_o;
  wire n7626_o;
  wire n7627_o;
  wire n7628_o;
  wire n7630_o;
  wire n7631_o;
  wire n7632_o;
  wire n7634_o;
  wire n7635_o;
  wire n7636_o;
  wire n7638_o;
  wire n7639_o;
  wire n7640_o;
  wire n7642_o;
  wire n7643_o;
  wire n7644_o;
  wire n7646_o;
  wire n7647_o;
  wire n7648_o;
  wire n7650_o;
  wire n7651_o;
  wire n7652_o;
  wire n7654_o;
  wire n7655_o;
  wire n7656_o;
  wire n7658_o;
  wire n7659_o;
  wire n7660_o;
  wire n7662_o;
  wire n7663_o;
  wire n7664_o;
  wire n7666_o;
  wire n7667_o;
  wire n7668_o;
  wire n7670_o;
  wire n7671_o;
  wire n7672_o;
  wire n7674_o;
  wire n7675_o;
  wire n7676_o;
  wire n7678_o;
  wire n7679_o;
  wire n7680_o;
  wire n7682_o;
  wire n7683_o;
  wire n7684_o;
  wire n7686_o;
  wire n7687_o;
  wire n7688_o;
  wire n7690_o;
  wire n7691_o;
  wire n7692_o;
  wire n7694_o;
  wire n7695_o;
  wire n7696_o;
  wire n7698_o;
  wire n7699_o;
  wire n7700_o;
  wire n7702_o;
  wire n7703_o;
  wire n7704_o;
  wire n7706_o;
  wire n7707_o;
  wire n7708_o;
  wire n7710_o;
  wire n7711_o;
  wire n7712_o;
  wire n7714_o;
  wire n7715_o;
  wire n7716_o;
  wire n7718_o;
  wire n7719_o;
  wire n7720_o;
  wire n7722_o;
  wire n7723_o;
  wire n7724_o;
  wire n7726_o;
  wire n7727_o;
  wire n7728_o;
  wire n7730_o;
  wire n7731_o;
  wire n7732_o;
  wire n7734_o;
  wire n7735_o;
  wire n7736_o;
  wire n7737_o;
  wire n7749_o;
  wire n7751_o;
  wire n7753_o;
  wire n7755_o;
  wire n7757_o;
  wire n7758_o;
  wire n7759_o;
  wire n7761_o;
  wire n7762_o;
  wire n7763_o;
  wire n7765_o;
  wire n7766_o;
  wire n7767_o;
  wire n7769_o;
  wire n7770_o;
  wire n7771_o;
  wire n7773_o;
  wire n7774_o;
  wire n7775_o;
  wire n7777_o;
  wire n7778_o;
  wire n7779_o;
  wire n7781_o;
  wire n7782_o;
  wire n7783_o;
  wire n7785_o;
  wire n7786_o;
  wire n7787_o;
  wire n7789_o;
  wire n7790_o;
  wire n7791_o;
  wire n7793_o;
  wire n7794_o;
  wire n7795_o;
  wire n7797_o;
  wire n7798_o;
  wire n7799_o;
  wire n7801_o;
  wire n7802_o;
  wire n7803_o;
  wire n7805_o;
  wire n7806_o;
  wire n7807_o;
  wire n7809_o;
  wire n7810_o;
  wire n7811_o;
  wire n7813_o;
  wire n7814_o;
  wire n7815_o;
  wire n7817_o;
  wire n7818_o;
  wire n7819_o;
  wire n7821_o;
  wire n7822_o;
  wire n7823_o;
  wire n7825_o;
  wire n7826_o;
  wire n7827_o;
  wire n7829_o;
  wire n7830_o;
  wire n7831_o;
  wire n7833_o;
  wire n7834_o;
  wire n7835_o;
  wire n7837_o;
  wire n7838_o;
  wire n7839_o;
  wire n7841_o;
  wire n7842_o;
  wire n7843_o;
  wire n7845_o;
  wire n7846_o;
  wire n7847_o;
  wire n7849_o;
  wire n7850_o;
  wire n7851_o;
  wire n7853_o;
  wire n7854_o;
  wire n7855_o;
  wire n7857_o;
  wire n7858_o;
  wire n7859_o;
  wire n7861_o;
  wire n7862_o;
  wire n7863_o;
  wire n7865_o;
  wire n7866_o;
  wire n7867_o;
  wire n7869_o;
  wire n7870_o;
  wire n7871_o;
  wire n7873_o;
  wire n7874_o;
  wire n7875_o;
  wire n7877_o;
  wire n7878_o;
  wire n7879_o;
  wire n7880_o;
  wire n7892_o;
  wire n7894_o;
  wire n7896_o;
  wire n7898_o;
  wire n7900_o;
  wire n7901_o;
  wire n7902_o;
  wire n7904_o;
  wire n7905_o;
  wire n7906_o;
  wire n7908_o;
  wire n7909_o;
  wire n7910_o;
  wire n7912_o;
  wire n7913_o;
  wire n7914_o;
  wire n7916_o;
  wire n7917_o;
  wire n7918_o;
  wire n7920_o;
  wire n7921_o;
  wire n7922_o;
  wire n7924_o;
  wire n7925_o;
  wire n7926_o;
  wire n7928_o;
  wire n7929_o;
  wire n7930_o;
  wire n7932_o;
  wire n7933_o;
  wire n7934_o;
  wire n7936_o;
  wire n7937_o;
  wire n7938_o;
  wire n7940_o;
  wire n7941_o;
  wire n7942_o;
  wire n7944_o;
  wire n7945_o;
  wire n7946_o;
  wire n7948_o;
  wire n7949_o;
  wire n7950_o;
  wire n7952_o;
  wire n7953_o;
  wire n7954_o;
  wire n7956_o;
  wire n7957_o;
  wire n7958_o;
  wire n7960_o;
  wire n7961_o;
  wire n7962_o;
  wire n7964_o;
  wire n7965_o;
  wire n7966_o;
  wire n7968_o;
  wire n7969_o;
  wire n7970_o;
  wire n7972_o;
  wire n7973_o;
  wire n7974_o;
  wire n7976_o;
  wire n7977_o;
  wire n7978_o;
  wire n7980_o;
  wire n7981_o;
  wire n7982_o;
  wire n7984_o;
  wire n7985_o;
  wire n7986_o;
  wire n7988_o;
  wire n7989_o;
  wire n7990_o;
  wire n7992_o;
  wire n7993_o;
  wire n7994_o;
  wire n7996_o;
  wire n7997_o;
  wire n7998_o;
  wire n8000_o;
  wire n8001_o;
  wire n8002_o;
  wire n8004_o;
  wire n8005_o;
  wire n8006_o;
  wire n8008_o;
  wire n8009_o;
  wire n8010_o;
  wire n8012_o;
  wire n8013_o;
  wire n8014_o;
  wire n8016_o;
  wire n8017_o;
  wire n8018_o;
  wire n8020_o;
  wire n8021_o;
  wire n8022_o;
  wire n8023_o;
  wire n8035_o;
  wire n8037_o;
  wire n8039_o;
  wire n8041_o;
  wire n8043_o;
  wire n8044_o;
  wire n8045_o;
  wire n8047_o;
  wire n8048_o;
  wire n8049_o;
  wire n8051_o;
  wire n8052_o;
  wire n8053_o;
  wire n8055_o;
  wire n8056_o;
  wire n8057_o;
  wire n8059_o;
  wire n8060_o;
  wire n8061_o;
  wire n8063_o;
  wire n8064_o;
  wire n8065_o;
  wire n8067_o;
  wire n8068_o;
  wire n8069_o;
  wire n8071_o;
  wire n8072_o;
  wire n8073_o;
  wire n8075_o;
  wire n8076_o;
  wire n8077_o;
  wire n8079_o;
  wire n8080_o;
  wire n8081_o;
  wire n8083_o;
  wire n8084_o;
  wire n8085_o;
  wire n8087_o;
  wire n8088_o;
  wire n8089_o;
  wire n8091_o;
  wire n8092_o;
  wire n8093_o;
  wire n8095_o;
  wire n8096_o;
  wire n8097_o;
  wire n8099_o;
  wire n8100_o;
  wire n8101_o;
  wire n8103_o;
  wire n8104_o;
  wire n8105_o;
  wire n8107_o;
  wire n8108_o;
  wire n8109_o;
  wire n8111_o;
  wire n8112_o;
  wire n8113_o;
  wire n8115_o;
  wire n8116_o;
  wire n8117_o;
  wire n8119_o;
  wire n8120_o;
  wire n8121_o;
  wire n8123_o;
  wire n8124_o;
  wire n8125_o;
  wire n8127_o;
  wire n8128_o;
  wire n8129_o;
  wire n8131_o;
  wire n8132_o;
  wire n8133_o;
  wire n8135_o;
  wire n8136_o;
  wire n8137_o;
  wire n8139_o;
  wire n8140_o;
  wire n8141_o;
  wire n8143_o;
  wire n8144_o;
  wire n8145_o;
  wire n8147_o;
  wire n8148_o;
  wire n8149_o;
  wire n8151_o;
  wire n8152_o;
  wire n8153_o;
  wire n8155_o;
  wire n8156_o;
  wire n8157_o;
  wire n8159_o;
  wire n8160_o;
  wire n8161_o;
  wire n8163_o;
  wire n8164_o;
  wire n8165_o;
  wire n8166_o;
  wire n8178_o;
  wire n8180_o;
  wire n8182_o;
  wire n8184_o;
  wire n8186_o;
  wire n8187_o;
  wire n8188_o;
  wire n8190_o;
  wire n8191_o;
  wire n8192_o;
  wire n8194_o;
  wire n8195_o;
  wire n8196_o;
  wire n8198_o;
  wire n8199_o;
  wire n8200_o;
  wire n8202_o;
  wire n8203_o;
  wire n8204_o;
  wire n8206_o;
  wire n8207_o;
  wire n8208_o;
  wire n8210_o;
  wire n8211_o;
  wire n8212_o;
  wire n8214_o;
  wire n8215_o;
  wire n8216_o;
  wire n8218_o;
  wire n8219_o;
  wire n8220_o;
  wire n8222_o;
  wire n8223_o;
  wire n8224_o;
  wire n8226_o;
  wire n8227_o;
  wire n8228_o;
  wire n8230_o;
  wire n8231_o;
  wire n8232_o;
  wire n8234_o;
  wire n8235_o;
  wire n8236_o;
  wire n8238_o;
  wire n8239_o;
  wire n8240_o;
  wire n8242_o;
  wire n8243_o;
  wire n8244_o;
  wire n8246_o;
  wire n8247_o;
  wire n8248_o;
  wire n8250_o;
  wire n8251_o;
  wire n8252_o;
  wire n8254_o;
  wire n8255_o;
  wire n8256_o;
  wire n8258_o;
  wire n8259_o;
  wire n8260_o;
  wire n8262_o;
  wire n8263_o;
  wire n8264_o;
  wire n8266_o;
  wire n8267_o;
  wire n8268_o;
  wire n8270_o;
  wire n8271_o;
  wire n8272_o;
  wire n8274_o;
  wire n8275_o;
  wire n8276_o;
  wire n8278_o;
  wire n8279_o;
  wire n8280_o;
  wire n8282_o;
  wire n8283_o;
  wire n8284_o;
  wire n8286_o;
  wire n8287_o;
  wire n8288_o;
  wire n8290_o;
  wire n8291_o;
  wire n8292_o;
  wire n8294_o;
  wire n8295_o;
  wire n8296_o;
  wire n8298_o;
  wire n8299_o;
  wire n8300_o;
  wire n8302_o;
  wire n8303_o;
  wire n8304_o;
  wire n8306_o;
  wire n8307_o;
  wire n8308_o;
  wire n8309_o;
  wire n8321_o;
  wire n8323_o;
  wire n8325_o;
  wire n8327_o;
  wire n8329_o;
  wire n8330_o;
  wire n8331_o;
  wire n8333_o;
  wire n8334_o;
  wire n8335_o;
  wire n8337_o;
  wire n8338_o;
  wire n8339_o;
  wire n8341_o;
  wire n8342_o;
  wire n8343_o;
  wire n8345_o;
  wire n8346_o;
  wire n8347_o;
  wire n8349_o;
  wire n8350_o;
  wire n8351_o;
  wire n8353_o;
  wire n8354_o;
  wire n8355_o;
  wire n8357_o;
  wire n8358_o;
  wire n8359_o;
  wire n8361_o;
  wire n8362_o;
  wire n8363_o;
  wire n8365_o;
  wire n8366_o;
  wire n8367_o;
  wire n8369_o;
  wire n8370_o;
  wire n8371_o;
  wire n8373_o;
  wire n8374_o;
  wire n8375_o;
  wire n8377_o;
  wire n8378_o;
  wire n8379_o;
  wire n8381_o;
  wire n8382_o;
  wire n8383_o;
  wire n8385_o;
  wire n8386_o;
  wire n8387_o;
  wire n8389_o;
  wire n8390_o;
  wire n8391_o;
  wire n8393_o;
  wire n8394_o;
  wire n8395_o;
  wire n8397_o;
  wire n8398_o;
  wire n8399_o;
  wire n8401_o;
  wire n8402_o;
  wire n8403_o;
  wire n8405_o;
  wire n8406_o;
  wire n8407_o;
  wire n8409_o;
  wire n8410_o;
  wire n8411_o;
  wire n8413_o;
  wire n8414_o;
  wire n8415_o;
  wire n8417_o;
  wire n8418_o;
  wire n8419_o;
  wire n8421_o;
  wire n8422_o;
  wire n8423_o;
  wire n8425_o;
  wire n8426_o;
  wire n8427_o;
  wire n8429_o;
  wire n8430_o;
  wire n8431_o;
  wire n8433_o;
  wire n8434_o;
  wire n8435_o;
  wire n8437_o;
  wire n8438_o;
  wire n8439_o;
  wire n8441_o;
  wire n8442_o;
  wire n8443_o;
  wire n8445_o;
  wire n8446_o;
  wire n8447_o;
  wire n8449_o;
  wire n8450_o;
  wire n8451_o;
  wire n8452_o;
  wire n8464_o;
  wire n8466_o;
  wire n8468_o;
  wire n8470_o;
  wire n8472_o;
  wire n8473_o;
  wire n8474_o;
  wire n8476_o;
  wire n8477_o;
  wire n8478_o;
  wire n8480_o;
  wire n8481_o;
  wire n8482_o;
  wire n8484_o;
  wire n8485_o;
  wire n8486_o;
  wire n8488_o;
  wire n8489_o;
  wire n8490_o;
  wire n8492_o;
  wire n8493_o;
  wire n8494_o;
  wire n8496_o;
  wire n8497_o;
  wire n8498_o;
  wire n8500_o;
  wire n8501_o;
  wire n8502_o;
  wire n8504_o;
  wire n8505_o;
  wire n8506_o;
  wire n8508_o;
  wire n8509_o;
  wire n8510_o;
  wire n8512_o;
  wire n8513_o;
  wire n8514_o;
  wire n8516_o;
  wire n8517_o;
  wire n8518_o;
  wire n8520_o;
  wire n8521_o;
  wire n8522_o;
  wire n8524_o;
  wire n8525_o;
  wire n8526_o;
  wire n8528_o;
  wire n8529_o;
  wire n8530_o;
  wire n8532_o;
  wire n8533_o;
  wire n8534_o;
  wire n8536_o;
  wire n8537_o;
  wire n8538_o;
  wire n8540_o;
  wire n8541_o;
  wire n8542_o;
  wire n8544_o;
  wire n8545_o;
  wire n8546_o;
  wire n8548_o;
  wire n8549_o;
  wire n8550_o;
  wire n8552_o;
  wire n8553_o;
  wire n8554_o;
  wire n8556_o;
  wire n8557_o;
  wire n8558_o;
  wire n8560_o;
  wire n8561_o;
  wire n8562_o;
  wire n8564_o;
  wire n8565_o;
  wire n8566_o;
  wire n8568_o;
  wire n8569_o;
  wire n8570_o;
  wire n8572_o;
  wire n8573_o;
  wire n8574_o;
  wire n8576_o;
  wire n8577_o;
  wire n8578_o;
  wire n8580_o;
  wire n8581_o;
  wire n8582_o;
  wire n8584_o;
  wire n8585_o;
  wire n8586_o;
  wire n8588_o;
  wire n8589_o;
  wire n8590_o;
  wire n8592_o;
  wire n8593_o;
  wire n8594_o;
  wire n8595_o;
  wire n8607_o;
  wire n8609_o;
  wire n8611_o;
  wire n8613_o;
  wire n8615_o;
  wire n8616_o;
  wire n8617_o;
  wire n8619_o;
  wire n8620_o;
  wire n8621_o;
  wire n8623_o;
  wire n8624_o;
  wire n8625_o;
  wire n8627_o;
  wire n8628_o;
  wire n8629_o;
  wire n8631_o;
  wire n8632_o;
  wire n8633_o;
  wire n8635_o;
  wire n8636_o;
  wire n8637_o;
  wire n8639_o;
  wire n8640_o;
  wire n8641_o;
  wire n8643_o;
  wire n8644_o;
  wire n8645_o;
  wire n8647_o;
  wire n8648_o;
  wire n8649_o;
  wire n8651_o;
  wire n8652_o;
  wire n8653_o;
  wire n8655_o;
  wire n8656_o;
  wire n8657_o;
  wire n8659_o;
  wire n8660_o;
  wire n8661_o;
  wire n8663_o;
  wire n8664_o;
  wire n8665_o;
  wire n8667_o;
  wire n8668_o;
  wire n8669_o;
  wire n8671_o;
  wire n8672_o;
  wire n8673_o;
  wire n8675_o;
  wire n8676_o;
  wire n8677_o;
  wire n8679_o;
  wire n8680_o;
  wire n8681_o;
  wire n8683_o;
  wire n8684_o;
  wire n8685_o;
  wire n8687_o;
  wire n8688_o;
  wire n8689_o;
  wire n8691_o;
  wire n8692_o;
  wire n8693_o;
  wire n8695_o;
  wire n8696_o;
  wire n8697_o;
  wire n8699_o;
  wire n8700_o;
  wire n8701_o;
  wire n8703_o;
  wire n8704_o;
  wire n8705_o;
  wire n8707_o;
  wire n8708_o;
  wire n8709_o;
  wire n8711_o;
  wire n8712_o;
  wire n8713_o;
  wire n8715_o;
  wire n8716_o;
  wire n8717_o;
  wire n8719_o;
  wire n8720_o;
  wire n8721_o;
  wire n8723_o;
  wire n8724_o;
  wire n8725_o;
  wire n8727_o;
  wire n8728_o;
  wire n8729_o;
  wire n8731_o;
  wire n8732_o;
  wire n8733_o;
  wire n8735_o;
  wire n8736_o;
  wire n8737_o;
  wire n8738_o;
  wire [3:0] n8739_o;
  wire [3:0] n8740_o;
  wire [1:0] n8741_o;
  wire [9:0] n8742_o;
  wire n8754_o;
  wire n8756_o;
  wire n8758_o;
  wire n8760_o;
  wire n8762_o;
  wire n8763_o;
  wire n8764_o;
  wire n8766_o;
  wire n8767_o;
  wire n8768_o;
  wire n8770_o;
  wire n8771_o;
  wire n8772_o;
  wire n8774_o;
  wire n8775_o;
  wire n8776_o;
  wire n8778_o;
  wire n8779_o;
  wire n8780_o;
  wire n8782_o;
  wire n8783_o;
  wire n8784_o;
  wire n8786_o;
  wire n8787_o;
  wire n8788_o;
  wire n8790_o;
  wire n8791_o;
  wire n8792_o;
  wire n8794_o;
  wire n8795_o;
  wire n8796_o;
  wire n8798_o;
  wire n8799_o;
  wire n8800_o;
  wire n8802_o;
  wire n8803_o;
  wire n8804_o;
  wire n8806_o;
  wire n8807_o;
  wire n8808_o;
  wire n8810_o;
  wire n8811_o;
  wire n8812_o;
  wire n8814_o;
  wire n8815_o;
  wire n8816_o;
  wire n8818_o;
  wire n8819_o;
  wire n8820_o;
  wire n8822_o;
  wire n8823_o;
  wire n8824_o;
  wire n8826_o;
  wire n8827_o;
  wire n8828_o;
  wire n8830_o;
  wire n8831_o;
  wire n8832_o;
  wire n8834_o;
  wire n8835_o;
  wire n8836_o;
  wire n8838_o;
  wire n8839_o;
  wire n8840_o;
  wire n8842_o;
  wire n8843_o;
  wire n8844_o;
  wire n8846_o;
  wire n8847_o;
  wire n8848_o;
  wire n8850_o;
  wire n8851_o;
  wire n8852_o;
  wire n8854_o;
  wire n8855_o;
  wire n8856_o;
  wire n8858_o;
  wire n8859_o;
  wire n8860_o;
  wire n8862_o;
  wire n8863_o;
  wire n8864_o;
  wire n8866_o;
  wire n8867_o;
  wire n8868_o;
  wire n8870_o;
  wire n8871_o;
  wire n8872_o;
  wire n8874_o;
  wire n8875_o;
  wire n8876_o;
  wire n8878_o;
  wire n8879_o;
  wire n8880_o;
  wire n8882_o;
  wire n8883_o;
  wire n8884_o;
  wire n8885_o;
  wire n8897_o;
  wire n8899_o;
  wire n8901_o;
  wire n8903_o;
  wire n8905_o;
  wire n8906_o;
  wire n8907_o;
  wire n8909_o;
  wire n8910_o;
  wire n8911_o;
  wire n8913_o;
  wire n8914_o;
  wire n8915_o;
  wire n8917_o;
  wire n8918_o;
  wire n8919_o;
  wire n8921_o;
  wire n8922_o;
  wire n8923_o;
  wire n8925_o;
  wire n8926_o;
  wire n8927_o;
  wire n8929_o;
  wire n8930_o;
  wire n8931_o;
  wire n8933_o;
  wire n8934_o;
  wire n8935_o;
  wire n8937_o;
  wire n8938_o;
  wire n8939_o;
  wire n8941_o;
  wire n8942_o;
  wire n8943_o;
  wire n8945_o;
  wire n8946_o;
  wire n8947_o;
  wire n8949_o;
  wire n8950_o;
  wire n8951_o;
  wire n8953_o;
  wire n8954_o;
  wire n8955_o;
  wire n8957_o;
  wire n8958_o;
  wire n8959_o;
  wire n8961_o;
  wire n8962_o;
  wire n8963_o;
  wire n8965_o;
  wire n8966_o;
  wire n8967_o;
  wire n8969_o;
  wire n8970_o;
  wire n8971_o;
  wire n8973_o;
  wire n8974_o;
  wire n8975_o;
  wire n8977_o;
  wire n8978_o;
  wire n8979_o;
  wire n8981_o;
  wire n8982_o;
  wire n8983_o;
  wire n8985_o;
  wire n8986_o;
  wire n8987_o;
  wire n8989_o;
  wire n8990_o;
  wire n8991_o;
  wire n8993_o;
  wire n8994_o;
  wire n8995_o;
  wire n8997_o;
  wire n8998_o;
  wire n8999_o;
  wire n9001_o;
  wire n9002_o;
  wire n9003_o;
  wire n9005_o;
  wire n9006_o;
  wire n9007_o;
  wire n9009_o;
  wire n9010_o;
  wire n9011_o;
  wire n9013_o;
  wire n9014_o;
  wire n9015_o;
  wire n9017_o;
  wire n9018_o;
  wire n9019_o;
  wire n9021_o;
  wire n9022_o;
  wire n9023_o;
  wire n9025_o;
  wire n9026_o;
  wire n9027_o;
  wire n9028_o;
  wire n9040_o;
  wire n9042_o;
  wire n9044_o;
  wire n9046_o;
  wire n9048_o;
  wire n9049_o;
  wire n9050_o;
  wire n9052_o;
  wire n9053_o;
  wire n9054_o;
  wire n9056_o;
  wire n9057_o;
  wire n9058_o;
  wire n9060_o;
  wire n9061_o;
  wire n9062_o;
  wire n9064_o;
  wire n9065_o;
  wire n9066_o;
  wire n9068_o;
  wire n9069_o;
  wire n9070_o;
  wire n9072_o;
  wire n9073_o;
  wire n9074_o;
  wire n9076_o;
  wire n9077_o;
  wire n9078_o;
  wire n9080_o;
  wire n9081_o;
  wire n9082_o;
  wire n9084_o;
  wire n9085_o;
  wire n9086_o;
  wire n9088_o;
  wire n9089_o;
  wire n9090_o;
  wire n9092_o;
  wire n9093_o;
  wire n9094_o;
  wire n9096_o;
  wire n9097_o;
  wire n9098_o;
  wire n9100_o;
  wire n9101_o;
  wire n9102_o;
  wire n9104_o;
  wire n9105_o;
  wire n9106_o;
  wire n9108_o;
  wire n9109_o;
  wire n9110_o;
  wire n9112_o;
  wire n9113_o;
  wire n9114_o;
  wire n9116_o;
  wire n9117_o;
  wire n9118_o;
  wire n9120_o;
  wire n9121_o;
  wire n9122_o;
  wire n9124_o;
  wire n9125_o;
  wire n9126_o;
  wire n9128_o;
  wire n9129_o;
  wire n9130_o;
  wire n9132_o;
  wire n9133_o;
  wire n9134_o;
  wire n9136_o;
  wire n9137_o;
  wire n9138_o;
  wire n9140_o;
  wire n9141_o;
  wire n9142_o;
  wire n9144_o;
  wire n9145_o;
  wire n9146_o;
  wire n9148_o;
  wire n9149_o;
  wire n9150_o;
  wire n9152_o;
  wire n9153_o;
  wire n9154_o;
  wire n9156_o;
  wire n9157_o;
  wire n9158_o;
  wire n9160_o;
  wire n9161_o;
  wire n9162_o;
  wire n9164_o;
  wire n9165_o;
  wire n9166_o;
  wire n9168_o;
  wire n9169_o;
  wire n9170_o;
  wire n9171_o;
  wire n9183_o;
  wire n9185_o;
  wire n9187_o;
  wire n9189_o;
  wire n9191_o;
  wire n9192_o;
  wire n9193_o;
  wire n9195_o;
  wire n9196_o;
  wire n9197_o;
  wire n9199_o;
  wire n9200_o;
  wire n9201_o;
  wire n9203_o;
  wire n9204_o;
  wire n9205_o;
  wire n9207_o;
  wire n9208_o;
  wire n9209_o;
  wire n9211_o;
  wire n9212_o;
  wire n9213_o;
  wire n9215_o;
  wire n9216_o;
  wire n9217_o;
  wire n9219_o;
  wire n9220_o;
  wire n9221_o;
  wire n9223_o;
  wire n9224_o;
  wire n9225_o;
  wire n9227_o;
  wire n9228_o;
  wire n9229_o;
  wire n9231_o;
  wire n9232_o;
  wire n9233_o;
  wire n9235_o;
  wire n9236_o;
  wire n9237_o;
  wire n9239_o;
  wire n9240_o;
  wire n9241_o;
  wire n9243_o;
  wire n9244_o;
  wire n9245_o;
  wire n9247_o;
  wire n9248_o;
  wire n9249_o;
  wire n9251_o;
  wire n9252_o;
  wire n9253_o;
  wire n9255_o;
  wire n9256_o;
  wire n9257_o;
  wire n9259_o;
  wire n9260_o;
  wire n9261_o;
  wire n9263_o;
  wire n9264_o;
  wire n9265_o;
  wire n9267_o;
  wire n9268_o;
  wire n9269_o;
  wire n9271_o;
  wire n9272_o;
  wire n9273_o;
  wire n9275_o;
  wire n9276_o;
  wire n9277_o;
  wire n9279_o;
  wire n9280_o;
  wire n9281_o;
  wire n9283_o;
  wire n9284_o;
  wire n9285_o;
  wire n9287_o;
  wire n9288_o;
  wire n9289_o;
  wire n9291_o;
  wire n9292_o;
  wire n9293_o;
  wire n9295_o;
  wire n9296_o;
  wire n9297_o;
  wire n9299_o;
  wire n9300_o;
  wire n9301_o;
  wire n9303_o;
  wire n9304_o;
  wire n9305_o;
  wire n9307_o;
  wire n9308_o;
  wire n9309_o;
  wire n9311_o;
  wire n9312_o;
  wire n9313_o;
  wire n9314_o;
  wire n9326_o;
  wire n9328_o;
  wire n9330_o;
  wire n9332_o;
  wire n9334_o;
  wire n9335_o;
  wire n9336_o;
  wire n9338_o;
  wire n9339_o;
  wire n9340_o;
  wire n9342_o;
  wire n9343_o;
  wire n9344_o;
  wire n9346_o;
  wire n9347_o;
  wire n9348_o;
  wire n9350_o;
  wire n9351_o;
  wire n9352_o;
  wire n9354_o;
  wire n9355_o;
  wire n9356_o;
  wire n9358_o;
  wire n9359_o;
  wire n9360_o;
  wire n9362_o;
  wire n9363_o;
  wire n9364_o;
  wire n9366_o;
  wire n9367_o;
  wire n9368_o;
  wire n9370_o;
  wire n9371_o;
  wire n9372_o;
  wire n9374_o;
  wire n9375_o;
  wire n9376_o;
  wire n9378_o;
  wire n9379_o;
  wire n9380_o;
  wire n9382_o;
  wire n9383_o;
  wire n9384_o;
  wire n9386_o;
  wire n9387_o;
  wire n9388_o;
  wire n9390_o;
  wire n9391_o;
  wire n9392_o;
  wire n9394_o;
  wire n9395_o;
  wire n9396_o;
  wire n9398_o;
  wire n9399_o;
  wire n9400_o;
  wire n9402_o;
  wire n9403_o;
  wire n9404_o;
  wire n9406_o;
  wire n9407_o;
  wire n9408_o;
  wire n9410_o;
  wire n9411_o;
  wire n9412_o;
  wire n9414_o;
  wire n9415_o;
  wire n9416_o;
  wire n9418_o;
  wire n9419_o;
  wire n9420_o;
  wire n9422_o;
  wire n9423_o;
  wire n9424_o;
  wire n9426_o;
  wire n9427_o;
  wire n9428_o;
  wire n9430_o;
  wire n9431_o;
  wire n9432_o;
  wire n9434_o;
  wire n9435_o;
  wire n9436_o;
  wire n9438_o;
  wire n9439_o;
  wire n9440_o;
  wire n9442_o;
  wire n9443_o;
  wire n9444_o;
  wire n9446_o;
  wire n9447_o;
  wire n9448_o;
  wire n9450_o;
  wire n9451_o;
  wire n9452_o;
  wire n9454_o;
  wire n9455_o;
  wire n9456_o;
  wire n9457_o;
  wire n9469_o;
  wire n9471_o;
  wire n9473_o;
  wire n9475_o;
  wire n9477_o;
  wire n9478_o;
  wire n9479_o;
  wire n9481_o;
  wire n9482_o;
  wire n9483_o;
  wire n9485_o;
  wire n9486_o;
  wire n9487_o;
  wire n9489_o;
  wire n9490_o;
  wire n9491_o;
  wire n9493_o;
  wire n9494_o;
  wire n9495_o;
  wire n9497_o;
  wire n9498_o;
  wire n9499_o;
  wire n9501_o;
  wire n9502_o;
  wire n9503_o;
  wire n9505_o;
  wire n9506_o;
  wire n9507_o;
  wire n9509_o;
  wire n9510_o;
  wire n9511_o;
  wire n9513_o;
  wire n9514_o;
  wire n9515_o;
  wire n9517_o;
  wire n9518_o;
  wire n9519_o;
  wire n9521_o;
  wire n9522_o;
  wire n9523_o;
  wire n9525_o;
  wire n9526_o;
  wire n9527_o;
  wire n9529_o;
  wire n9530_o;
  wire n9531_o;
  wire n9533_o;
  wire n9534_o;
  wire n9535_o;
  wire n9537_o;
  wire n9538_o;
  wire n9539_o;
  wire n9541_o;
  wire n9542_o;
  wire n9543_o;
  wire n9545_o;
  wire n9546_o;
  wire n9547_o;
  wire n9549_o;
  wire n9550_o;
  wire n9551_o;
  wire n9553_o;
  wire n9554_o;
  wire n9555_o;
  wire n9557_o;
  wire n9558_o;
  wire n9559_o;
  wire n9561_o;
  wire n9562_o;
  wire n9563_o;
  wire n9565_o;
  wire n9566_o;
  wire n9567_o;
  wire n9569_o;
  wire n9570_o;
  wire n9571_o;
  wire n9573_o;
  wire n9574_o;
  wire n9575_o;
  wire n9577_o;
  wire n9578_o;
  wire n9579_o;
  wire n9581_o;
  wire n9582_o;
  wire n9583_o;
  wire n9585_o;
  wire n9586_o;
  wire n9587_o;
  wire n9589_o;
  wire n9590_o;
  wire n9591_o;
  wire n9593_o;
  wire n9594_o;
  wire n9595_o;
  wire n9597_o;
  wire n9598_o;
  wire n9599_o;
  wire n9600_o;
  wire n9612_o;
  wire n9614_o;
  wire n9616_o;
  wire n9618_o;
  wire n9620_o;
  wire n9621_o;
  wire n9622_o;
  wire n9624_o;
  wire n9625_o;
  wire n9626_o;
  wire n9628_o;
  wire n9629_o;
  wire n9630_o;
  wire n9632_o;
  wire n9633_o;
  wire n9634_o;
  wire n9636_o;
  wire n9637_o;
  wire n9638_o;
  wire n9640_o;
  wire n9641_o;
  wire n9642_o;
  wire n9644_o;
  wire n9645_o;
  wire n9646_o;
  wire n9648_o;
  wire n9649_o;
  wire n9650_o;
  wire n9652_o;
  wire n9653_o;
  wire n9654_o;
  wire n9656_o;
  wire n9657_o;
  wire n9658_o;
  wire n9660_o;
  wire n9661_o;
  wire n9662_o;
  wire n9664_o;
  wire n9665_o;
  wire n9666_o;
  wire n9668_o;
  wire n9669_o;
  wire n9670_o;
  wire n9672_o;
  wire n9673_o;
  wire n9674_o;
  wire n9676_o;
  wire n9677_o;
  wire n9678_o;
  wire n9680_o;
  wire n9681_o;
  wire n9682_o;
  wire n9684_o;
  wire n9685_o;
  wire n9686_o;
  wire n9688_o;
  wire n9689_o;
  wire n9690_o;
  wire n9692_o;
  wire n9693_o;
  wire n9694_o;
  wire n9696_o;
  wire n9697_o;
  wire n9698_o;
  wire n9700_o;
  wire n9701_o;
  wire n9702_o;
  wire n9704_o;
  wire n9705_o;
  wire n9706_o;
  wire n9708_o;
  wire n9709_o;
  wire n9710_o;
  wire n9712_o;
  wire n9713_o;
  wire n9714_o;
  wire n9716_o;
  wire n9717_o;
  wire n9718_o;
  wire n9720_o;
  wire n9721_o;
  wire n9722_o;
  wire n9724_o;
  wire n9725_o;
  wire n9726_o;
  wire n9728_o;
  wire n9729_o;
  wire n9730_o;
  wire n9732_o;
  wire n9733_o;
  wire n9734_o;
  wire n9736_o;
  wire n9737_o;
  wire n9738_o;
  wire n9740_o;
  wire n9741_o;
  wire n9742_o;
  wire n9743_o;
  wire n9755_o;
  wire n9757_o;
  wire n9759_o;
  wire n9761_o;
  wire n9763_o;
  wire n9764_o;
  wire n9765_o;
  wire n9767_o;
  wire n9768_o;
  wire n9769_o;
  wire n9771_o;
  wire n9772_o;
  wire n9773_o;
  wire n9775_o;
  wire n9776_o;
  wire n9777_o;
  wire n9779_o;
  wire n9780_o;
  wire n9781_o;
  wire n9783_o;
  wire n9784_o;
  wire n9785_o;
  wire n9787_o;
  wire n9788_o;
  wire n9789_o;
  wire n9791_o;
  wire n9792_o;
  wire n9793_o;
  wire n9795_o;
  wire n9796_o;
  wire n9797_o;
  wire n9799_o;
  wire n9800_o;
  wire n9801_o;
  wire n9803_o;
  wire n9804_o;
  wire n9805_o;
  wire n9807_o;
  wire n9808_o;
  wire n9809_o;
  wire n9811_o;
  wire n9812_o;
  wire n9813_o;
  wire n9815_o;
  wire n9816_o;
  wire n9817_o;
  wire n9819_o;
  wire n9820_o;
  wire n9821_o;
  wire n9823_o;
  wire n9824_o;
  wire n9825_o;
  wire n9827_o;
  wire n9828_o;
  wire n9829_o;
  wire n9831_o;
  wire n9832_o;
  wire n9833_o;
  wire n9835_o;
  wire n9836_o;
  wire n9837_o;
  wire n9839_o;
  wire n9840_o;
  wire n9841_o;
  wire n9843_o;
  wire n9844_o;
  wire n9845_o;
  wire n9847_o;
  wire n9848_o;
  wire n9849_o;
  wire n9851_o;
  wire n9852_o;
  wire n9853_o;
  wire n9855_o;
  wire n9856_o;
  wire n9857_o;
  wire n9859_o;
  wire n9860_o;
  wire n9861_o;
  wire n9863_o;
  wire n9864_o;
  wire n9865_o;
  wire n9867_o;
  wire n9868_o;
  wire n9869_o;
  wire n9871_o;
  wire n9872_o;
  wire n9873_o;
  wire n9875_o;
  wire n9876_o;
  wire n9877_o;
  wire n9879_o;
  wire n9880_o;
  wire n9881_o;
  wire n9883_o;
  wire n9884_o;
  wire n9885_o;
  wire n9886_o;
  wire n9898_o;
  wire n9900_o;
  wire n9902_o;
  wire n9904_o;
  wire n9906_o;
  wire n9907_o;
  wire n9908_o;
  wire n9910_o;
  wire n9911_o;
  wire n9912_o;
  wire n9914_o;
  wire n9915_o;
  wire n9916_o;
  wire n9918_o;
  wire n9919_o;
  wire n9920_o;
  wire n9922_o;
  wire n9923_o;
  wire n9924_o;
  wire n9926_o;
  wire n9927_o;
  wire n9928_o;
  wire n9930_o;
  wire n9931_o;
  wire n9932_o;
  wire n9934_o;
  wire n9935_o;
  wire n9936_o;
  wire n9938_o;
  wire n9939_o;
  wire n9940_o;
  wire n9942_o;
  wire n9943_o;
  wire n9944_o;
  wire n9946_o;
  wire n9947_o;
  wire n9948_o;
  wire n9950_o;
  wire n9951_o;
  wire n9952_o;
  wire n9954_o;
  wire n9955_o;
  wire n9956_o;
  wire n9958_o;
  wire n9959_o;
  wire n9960_o;
  wire n9962_o;
  wire n9963_o;
  wire n9964_o;
  wire n9966_o;
  wire n9967_o;
  wire n9968_o;
  wire n9970_o;
  wire n9971_o;
  wire n9972_o;
  wire n9974_o;
  wire n9975_o;
  wire n9976_o;
  wire n9978_o;
  wire n9979_o;
  wire n9980_o;
  wire n9982_o;
  wire n9983_o;
  wire n9984_o;
  wire n9986_o;
  wire n9987_o;
  wire n9988_o;
  wire n9990_o;
  wire n9991_o;
  wire n9992_o;
  wire n9994_o;
  wire n9995_o;
  wire n9996_o;
  wire n9998_o;
  wire n9999_o;
  wire n10000_o;
  wire n10002_o;
  wire n10003_o;
  wire n10004_o;
  wire n10006_o;
  wire n10007_o;
  wire n10008_o;
  wire n10010_o;
  wire n10011_o;
  wire n10012_o;
  wire n10014_o;
  wire n10015_o;
  wire n10016_o;
  wire n10018_o;
  wire n10019_o;
  wire n10020_o;
  wire n10022_o;
  wire n10023_o;
  wire n10024_o;
  wire n10026_o;
  wire n10027_o;
  wire n10028_o;
  wire n10029_o;
  wire n10041_o;
  wire n10043_o;
  wire n10045_o;
  wire n10047_o;
  wire n10049_o;
  wire n10050_o;
  wire n10051_o;
  wire n10053_o;
  wire n10054_o;
  wire n10055_o;
  wire n10057_o;
  wire n10058_o;
  wire n10059_o;
  wire n10061_o;
  wire n10062_o;
  wire n10063_o;
  wire n10065_o;
  wire n10066_o;
  wire n10067_o;
  wire n10069_o;
  wire n10070_o;
  wire n10071_o;
  wire n10073_o;
  wire n10074_o;
  wire n10075_o;
  wire n10077_o;
  wire n10078_o;
  wire n10079_o;
  wire n10081_o;
  wire n10082_o;
  wire n10083_o;
  wire n10085_o;
  wire n10086_o;
  wire n10087_o;
  wire n10089_o;
  wire n10090_o;
  wire n10091_o;
  wire n10093_o;
  wire n10094_o;
  wire n10095_o;
  wire n10097_o;
  wire n10098_o;
  wire n10099_o;
  wire n10101_o;
  wire n10102_o;
  wire n10103_o;
  wire n10105_o;
  wire n10106_o;
  wire n10107_o;
  wire n10109_o;
  wire n10110_o;
  wire n10111_o;
  wire n10113_o;
  wire n10114_o;
  wire n10115_o;
  wire n10117_o;
  wire n10118_o;
  wire n10119_o;
  wire n10121_o;
  wire n10122_o;
  wire n10123_o;
  wire n10125_o;
  wire n10126_o;
  wire n10127_o;
  wire n10129_o;
  wire n10130_o;
  wire n10131_o;
  wire n10133_o;
  wire n10134_o;
  wire n10135_o;
  wire n10137_o;
  wire n10138_o;
  wire n10139_o;
  wire n10141_o;
  wire n10142_o;
  wire n10143_o;
  wire n10145_o;
  wire n10146_o;
  wire n10147_o;
  wire n10149_o;
  wire n10150_o;
  wire n10151_o;
  wire n10153_o;
  wire n10154_o;
  wire n10155_o;
  wire n10157_o;
  wire n10158_o;
  wire n10159_o;
  wire n10161_o;
  wire n10162_o;
  wire n10163_o;
  wire n10165_o;
  wire n10166_o;
  wire n10167_o;
  wire n10169_o;
  wire n10170_o;
  wire n10171_o;
  wire n10172_o;
  wire [3:0] n10173_o;
  wire [3:0] n10174_o;
  wire [1:0] n10175_o;
  wire [9:0] n10176_o;
  wire n10188_o;
  wire n10190_o;
  wire n10192_o;
  wire n10194_o;
  wire n10196_o;
  wire n10197_o;
  wire n10198_o;
  wire n10200_o;
  wire n10201_o;
  wire n10202_o;
  wire n10204_o;
  wire n10205_o;
  wire n10206_o;
  wire n10208_o;
  wire n10209_o;
  wire n10210_o;
  wire n10212_o;
  wire n10213_o;
  wire n10214_o;
  wire n10216_o;
  wire n10217_o;
  wire n10218_o;
  wire n10220_o;
  wire n10221_o;
  wire n10222_o;
  wire n10224_o;
  wire n10225_o;
  wire n10226_o;
  wire n10228_o;
  wire n10229_o;
  wire n10230_o;
  wire n10232_o;
  wire n10233_o;
  wire n10234_o;
  wire n10236_o;
  wire n10237_o;
  wire n10238_o;
  wire n10240_o;
  wire n10241_o;
  wire n10242_o;
  wire n10244_o;
  wire n10245_o;
  wire n10246_o;
  wire n10248_o;
  wire n10249_o;
  wire n10250_o;
  wire n10252_o;
  wire n10253_o;
  wire n10254_o;
  wire n10256_o;
  wire n10257_o;
  wire n10258_o;
  wire n10260_o;
  wire n10261_o;
  wire n10262_o;
  wire n10264_o;
  wire n10265_o;
  wire n10266_o;
  wire n10268_o;
  wire n10269_o;
  wire n10270_o;
  wire n10272_o;
  wire n10273_o;
  wire n10274_o;
  wire n10276_o;
  wire n10277_o;
  wire n10278_o;
  wire n10280_o;
  wire n10281_o;
  wire n10282_o;
  wire n10284_o;
  wire n10285_o;
  wire n10286_o;
  wire n10288_o;
  wire n10289_o;
  wire n10290_o;
  wire n10292_o;
  wire n10293_o;
  wire n10294_o;
  wire n10296_o;
  wire n10297_o;
  wire n10298_o;
  wire n10300_o;
  wire n10301_o;
  wire n10302_o;
  wire n10304_o;
  wire n10305_o;
  wire n10306_o;
  wire n10308_o;
  wire n10309_o;
  wire n10310_o;
  wire n10312_o;
  wire n10313_o;
  wire n10314_o;
  wire n10316_o;
  wire n10317_o;
  wire n10318_o;
  wire n10319_o;
  wire n10331_o;
  wire n10333_o;
  wire n10335_o;
  wire n10337_o;
  wire n10339_o;
  wire n10340_o;
  wire n10341_o;
  wire n10343_o;
  wire n10344_o;
  wire n10345_o;
  wire n10347_o;
  wire n10348_o;
  wire n10349_o;
  wire n10351_o;
  wire n10352_o;
  wire n10353_o;
  wire n10355_o;
  wire n10356_o;
  wire n10357_o;
  wire n10359_o;
  wire n10360_o;
  wire n10361_o;
  wire n10363_o;
  wire n10364_o;
  wire n10365_o;
  wire n10367_o;
  wire n10368_o;
  wire n10369_o;
  wire n10371_o;
  wire n10372_o;
  wire n10373_o;
  wire n10375_o;
  wire n10376_o;
  wire n10377_o;
  wire n10379_o;
  wire n10380_o;
  wire n10381_o;
  wire n10383_o;
  wire n10384_o;
  wire n10385_o;
  wire n10387_o;
  wire n10388_o;
  wire n10389_o;
  wire n10391_o;
  wire n10392_o;
  wire n10393_o;
  wire n10395_o;
  wire n10396_o;
  wire n10397_o;
  wire n10399_o;
  wire n10400_o;
  wire n10401_o;
  wire n10403_o;
  wire n10404_o;
  wire n10405_o;
  wire n10407_o;
  wire n10408_o;
  wire n10409_o;
  wire n10411_o;
  wire n10412_o;
  wire n10413_o;
  wire n10415_o;
  wire n10416_o;
  wire n10417_o;
  wire n10419_o;
  wire n10420_o;
  wire n10421_o;
  wire n10423_o;
  wire n10424_o;
  wire n10425_o;
  wire n10427_o;
  wire n10428_o;
  wire n10429_o;
  wire n10431_o;
  wire n10432_o;
  wire n10433_o;
  wire n10435_o;
  wire n10436_o;
  wire n10437_o;
  wire n10439_o;
  wire n10440_o;
  wire n10441_o;
  wire n10443_o;
  wire n10444_o;
  wire n10445_o;
  wire n10447_o;
  wire n10448_o;
  wire n10449_o;
  wire n10451_o;
  wire n10452_o;
  wire n10453_o;
  wire n10455_o;
  wire n10456_o;
  wire n10457_o;
  wire n10459_o;
  wire n10460_o;
  wire n10461_o;
  wire n10462_o;
  wire n10474_o;
  wire n10476_o;
  wire n10478_o;
  wire n10480_o;
  wire n10482_o;
  wire n10483_o;
  wire n10484_o;
  wire n10486_o;
  wire n10487_o;
  wire n10488_o;
  wire n10490_o;
  wire n10491_o;
  wire n10492_o;
  wire n10494_o;
  wire n10495_o;
  wire n10496_o;
  wire n10498_o;
  wire n10499_o;
  wire n10500_o;
  wire n10502_o;
  wire n10503_o;
  wire n10504_o;
  wire n10506_o;
  wire n10507_o;
  wire n10508_o;
  wire n10510_o;
  wire n10511_o;
  wire n10512_o;
  wire n10514_o;
  wire n10515_o;
  wire n10516_o;
  wire n10518_o;
  wire n10519_o;
  wire n10520_o;
  wire n10522_o;
  wire n10523_o;
  wire n10524_o;
  wire n10526_o;
  wire n10527_o;
  wire n10528_o;
  wire n10530_o;
  wire n10531_o;
  wire n10532_o;
  wire n10534_o;
  wire n10535_o;
  wire n10536_o;
  wire n10538_o;
  wire n10539_o;
  wire n10540_o;
  wire n10542_o;
  wire n10543_o;
  wire n10544_o;
  wire n10546_o;
  wire n10547_o;
  wire n10548_o;
  wire n10550_o;
  wire n10551_o;
  wire n10552_o;
  wire n10554_o;
  wire n10555_o;
  wire n10556_o;
  wire n10558_o;
  wire n10559_o;
  wire n10560_o;
  wire n10562_o;
  wire n10563_o;
  wire n10564_o;
  wire n10566_o;
  wire n10567_o;
  wire n10568_o;
  wire n10570_o;
  wire n10571_o;
  wire n10572_o;
  wire n10574_o;
  wire n10575_o;
  wire n10576_o;
  wire n10578_o;
  wire n10579_o;
  wire n10580_o;
  wire n10582_o;
  wire n10583_o;
  wire n10584_o;
  wire n10586_o;
  wire n10587_o;
  wire n10588_o;
  wire n10590_o;
  wire n10591_o;
  wire n10592_o;
  wire n10594_o;
  wire n10595_o;
  wire n10596_o;
  wire n10598_o;
  wire n10599_o;
  wire n10600_o;
  wire n10602_o;
  wire n10603_o;
  wire n10604_o;
  wire n10605_o;
  wire n10617_o;
  wire n10619_o;
  wire n10621_o;
  wire n10623_o;
  wire n10625_o;
  wire n10626_o;
  wire n10627_o;
  wire n10629_o;
  wire n10630_o;
  wire n10631_o;
  wire n10633_o;
  wire n10634_o;
  wire n10635_o;
  wire n10637_o;
  wire n10638_o;
  wire n10639_o;
  wire n10641_o;
  wire n10642_o;
  wire n10643_o;
  wire n10645_o;
  wire n10646_o;
  wire n10647_o;
  wire n10649_o;
  wire n10650_o;
  wire n10651_o;
  wire n10653_o;
  wire n10654_o;
  wire n10655_o;
  wire n10657_o;
  wire n10658_o;
  wire n10659_o;
  wire n10661_o;
  wire n10662_o;
  wire n10663_o;
  wire n10665_o;
  wire n10666_o;
  wire n10667_o;
  wire n10669_o;
  wire n10670_o;
  wire n10671_o;
  wire n10673_o;
  wire n10674_o;
  wire n10675_o;
  wire n10677_o;
  wire n10678_o;
  wire n10679_o;
  wire n10681_o;
  wire n10682_o;
  wire n10683_o;
  wire n10685_o;
  wire n10686_o;
  wire n10687_o;
  wire n10689_o;
  wire n10690_o;
  wire n10691_o;
  wire n10693_o;
  wire n10694_o;
  wire n10695_o;
  wire n10697_o;
  wire n10698_o;
  wire n10699_o;
  wire n10701_o;
  wire n10702_o;
  wire n10703_o;
  wire n10705_o;
  wire n10706_o;
  wire n10707_o;
  wire n10709_o;
  wire n10710_o;
  wire n10711_o;
  wire n10713_o;
  wire n10714_o;
  wire n10715_o;
  wire n10717_o;
  wire n10718_o;
  wire n10719_o;
  wire n10721_o;
  wire n10722_o;
  wire n10723_o;
  wire n10725_o;
  wire n10726_o;
  wire n10727_o;
  wire n10729_o;
  wire n10730_o;
  wire n10731_o;
  wire n10733_o;
  wire n10734_o;
  wire n10735_o;
  wire n10737_o;
  wire n10738_o;
  wire n10739_o;
  wire n10741_o;
  wire n10742_o;
  wire n10743_o;
  wire n10745_o;
  wire n10746_o;
  wire n10747_o;
  wire n10748_o;
  wire n10760_o;
  wire n10762_o;
  wire n10764_o;
  wire n10766_o;
  wire n10768_o;
  wire n10769_o;
  wire n10770_o;
  wire n10772_o;
  wire n10773_o;
  wire n10774_o;
  wire n10776_o;
  wire n10777_o;
  wire n10778_o;
  wire n10780_o;
  wire n10781_o;
  wire n10782_o;
  wire n10784_o;
  wire n10785_o;
  wire n10786_o;
  wire n10788_o;
  wire n10789_o;
  wire n10790_o;
  wire n10792_o;
  wire n10793_o;
  wire n10794_o;
  wire n10796_o;
  wire n10797_o;
  wire n10798_o;
  wire n10800_o;
  wire n10801_o;
  wire n10802_o;
  wire n10804_o;
  wire n10805_o;
  wire n10806_o;
  wire n10808_o;
  wire n10809_o;
  wire n10810_o;
  wire n10812_o;
  wire n10813_o;
  wire n10814_o;
  wire n10816_o;
  wire n10817_o;
  wire n10818_o;
  wire n10820_o;
  wire n10821_o;
  wire n10822_o;
  wire n10824_o;
  wire n10825_o;
  wire n10826_o;
  wire n10828_o;
  wire n10829_o;
  wire n10830_o;
  wire n10832_o;
  wire n10833_o;
  wire n10834_o;
  wire n10836_o;
  wire n10837_o;
  wire n10838_o;
  wire n10840_o;
  wire n10841_o;
  wire n10842_o;
  wire n10844_o;
  wire n10845_o;
  wire n10846_o;
  wire n10848_o;
  wire n10849_o;
  wire n10850_o;
  wire n10852_o;
  wire n10853_o;
  wire n10854_o;
  wire n10856_o;
  wire n10857_o;
  wire n10858_o;
  wire n10860_o;
  wire n10861_o;
  wire n10862_o;
  wire n10864_o;
  wire n10865_o;
  wire n10866_o;
  wire n10868_o;
  wire n10869_o;
  wire n10870_o;
  wire n10872_o;
  wire n10873_o;
  wire n10874_o;
  wire n10876_o;
  wire n10877_o;
  wire n10878_o;
  wire n10880_o;
  wire n10881_o;
  wire n10882_o;
  wire n10884_o;
  wire n10885_o;
  wire n10886_o;
  wire n10888_o;
  wire n10889_o;
  wire n10890_o;
  wire n10891_o;
  wire n10903_o;
  wire n10905_o;
  wire n10907_o;
  wire n10909_o;
  wire n10911_o;
  wire n10912_o;
  wire n10913_o;
  wire n10915_o;
  wire n10916_o;
  wire n10917_o;
  wire n10919_o;
  wire n10920_o;
  wire n10921_o;
  wire n10923_o;
  wire n10924_o;
  wire n10925_o;
  wire n10927_o;
  wire n10928_o;
  wire n10929_o;
  wire n10931_o;
  wire n10932_o;
  wire n10933_o;
  wire n10935_o;
  wire n10936_o;
  wire n10937_o;
  wire n10939_o;
  wire n10940_o;
  wire n10941_o;
  wire n10943_o;
  wire n10944_o;
  wire n10945_o;
  wire n10947_o;
  wire n10948_o;
  wire n10949_o;
  wire n10951_o;
  wire n10952_o;
  wire n10953_o;
  wire n10955_o;
  wire n10956_o;
  wire n10957_o;
  wire n10959_o;
  wire n10960_o;
  wire n10961_o;
  wire n10963_o;
  wire n10964_o;
  wire n10965_o;
  wire n10967_o;
  wire n10968_o;
  wire n10969_o;
  wire n10971_o;
  wire n10972_o;
  wire n10973_o;
  wire n10975_o;
  wire n10976_o;
  wire n10977_o;
  wire n10979_o;
  wire n10980_o;
  wire n10981_o;
  wire n10983_o;
  wire n10984_o;
  wire n10985_o;
  wire n10987_o;
  wire n10988_o;
  wire n10989_o;
  wire n10991_o;
  wire n10992_o;
  wire n10993_o;
  wire n10995_o;
  wire n10996_o;
  wire n10997_o;
  wire n10999_o;
  wire n11000_o;
  wire n11001_o;
  wire n11003_o;
  wire n11004_o;
  wire n11005_o;
  wire n11007_o;
  wire n11008_o;
  wire n11009_o;
  wire n11011_o;
  wire n11012_o;
  wire n11013_o;
  wire n11015_o;
  wire n11016_o;
  wire n11017_o;
  wire n11019_o;
  wire n11020_o;
  wire n11021_o;
  wire n11023_o;
  wire n11024_o;
  wire n11025_o;
  wire n11027_o;
  wire n11028_o;
  wire n11029_o;
  wire n11031_o;
  wire n11032_o;
  wire n11033_o;
  wire n11034_o;
  wire n11046_o;
  wire n11048_o;
  wire n11050_o;
  wire n11052_o;
  wire n11054_o;
  wire n11055_o;
  wire n11056_o;
  wire n11058_o;
  wire n11059_o;
  wire n11060_o;
  wire n11062_o;
  wire n11063_o;
  wire n11064_o;
  wire n11066_o;
  wire n11067_o;
  wire n11068_o;
  wire n11070_o;
  wire n11071_o;
  wire n11072_o;
  wire n11074_o;
  wire n11075_o;
  wire n11076_o;
  wire n11078_o;
  wire n11079_o;
  wire n11080_o;
  wire n11082_o;
  wire n11083_o;
  wire n11084_o;
  wire n11086_o;
  wire n11087_o;
  wire n11088_o;
  wire n11090_o;
  wire n11091_o;
  wire n11092_o;
  wire n11094_o;
  wire n11095_o;
  wire n11096_o;
  wire n11098_o;
  wire n11099_o;
  wire n11100_o;
  wire n11102_o;
  wire n11103_o;
  wire n11104_o;
  wire n11106_o;
  wire n11107_o;
  wire n11108_o;
  wire n11110_o;
  wire n11111_o;
  wire n11112_o;
  wire n11114_o;
  wire n11115_o;
  wire n11116_o;
  wire n11118_o;
  wire n11119_o;
  wire n11120_o;
  wire n11122_o;
  wire n11123_o;
  wire n11124_o;
  wire n11126_o;
  wire n11127_o;
  wire n11128_o;
  wire n11130_o;
  wire n11131_o;
  wire n11132_o;
  wire n11134_o;
  wire n11135_o;
  wire n11136_o;
  wire n11138_o;
  wire n11139_o;
  wire n11140_o;
  wire n11142_o;
  wire n11143_o;
  wire n11144_o;
  wire n11146_o;
  wire n11147_o;
  wire n11148_o;
  wire n11150_o;
  wire n11151_o;
  wire n11152_o;
  wire n11154_o;
  wire n11155_o;
  wire n11156_o;
  wire n11158_o;
  wire n11159_o;
  wire n11160_o;
  wire n11162_o;
  wire n11163_o;
  wire n11164_o;
  wire n11166_o;
  wire n11167_o;
  wire n11168_o;
  wire n11170_o;
  wire n11171_o;
  wire n11172_o;
  wire n11174_o;
  wire n11175_o;
  wire n11176_o;
  wire n11177_o;
  wire [3:0] n11181_o;
  wire [3:0] n11182_o;
  wire [1:0] n11183_o;
  wire [9:0] n11184_o;
  wire n11196_o;
  wire n11198_o;
  wire n11200_o;
  wire n11202_o;
  wire n11204_o;
  wire n11205_o;
  wire n11206_o;
  wire n11208_o;
  wire n11209_o;
  wire n11210_o;
  wire n11212_o;
  wire n11213_o;
  wire n11214_o;
  wire n11216_o;
  wire n11217_o;
  wire n11218_o;
  wire n11220_o;
  wire n11221_o;
  wire n11222_o;
  wire n11224_o;
  wire n11225_o;
  wire n11226_o;
  wire n11228_o;
  wire n11229_o;
  wire n11230_o;
  wire n11232_o;
  wire n11233_o;
  wire n11234_o;
  wire n11236_o;
  wire n11237_o;
  wire n11238_o;
  wire n11240_o;
  wire n11241_o;
  wire n11242_o;
  wire n11244_o;
  wire n11245_o;
  wire n11246_o;
  wire n11248_o;
  wire n11249_o;
  wire n11250_o;
  wire n11252_o;
  wire n11253_o;
  wire n11254_o;
  wire n11256_o;
  wire n11257_o;
  wire n11258_o;
  wire n11260_o;
  wire n11261_o;
  wire n11262_o;
  wire n11264_o;
  wire n11265_o;
  wire n11266_o;
  wire n11268_o;
  wire n11269_o;
  wire n11270_o;
  wire n11272_o;
  wire n11273_o;
  wire n11274_o;
  wire n11276_o;
  wire n11277_o;
  wire n11278_o;
  wire n11280_o;
  wire n11281_o;
  wire n11282_o;
  wire n11284_o;
  wire n11285_o;
  wire n11286_o;
  wire n11288_o;
  wire n11289_o;
  wire n11290_o;
  wire n11292_o;
  wire n11293_o;
  wire n11294_o;
  wire n11296_o;
  wire n11297_o;
  wire n11298_o;
  wire n11300_o;
  wire n11301_o;
  wire n11302_o;
  wire n11304_o;
  wire n11305_o;
  wire n11306_o;
  wire n11308_o;
  wire n11309_o;
  wire n11310_o;
  wire n11312_o;
  wire n11313_o;
  wire n11314_o;
  wire n11316_o;
  wire n11317_o;
  wire n11318_o;
  wire n11320_o;
  wire n11321_o;
  wire n11322_o;
  wire n11324_o;
  wire n11325_o;
  wire n11326_o;
  wire n11327_o;
  wire n11339_o;
  wire n11341_o;
  wire n11343_o;
  wire n11345_o;
  wire n11347_o;
  wire n11348_o;
  wire n11349_o;
  wire n11351_o;
  wire n11352_o;
  wire n11353_o;
  wire n11355_o;
  wire n11356_o;
  wire n11357_o;
  wire n11359_o;
  wire n11360_o;
  wire n11361_o;
  wire n11363_o;
  wire n11364_o;
  wire n11365_o;
  wire n11367_o;
  wire n11368_o;
  wire n11369_o;
  wire n11371_o;
  wire n11372_o;
  wire n11373_o;
  wire n11375_o;
  wire n11376_o;
  wire n11377_o;
  wire n11379_o;
  wire n11380_o;
  wire n11381_o;
  wire n11383_o;
  wire n11384_o;
  wire n11385_o;
  wire n11387_o;
  wire n11388_o;
  wire n11389_o;
  wire n11391_o;
  wire n11392_o;
  wire n11393_o;
  wire n11395_o;
  wire n11396_o;
  wire n11397_o;
  wire n11399_o;
  wire n11400_o;
  wire n11401_o;
  wire n11403_o;
  wire n11404_o;
  wire n11405_o;
  wire n11407_o;
  wire n11408_o;
  wire n11409_o;
  wire n11411_o;
  wire n11412_o;
  wire n11413_o;
  wire n11415_o;
  wire n11416_o;
  wire n11417_o;
  wire n11419_o;
  wire n11420_o;
  wire n11421_o;
  wire n11423_o;
  wire n11424_o;
  wire n11425_o;
  wire n11427_o;
  wire n11428_o;
  wire n11429_o;
  wire n11431_o;
  wire n11432_o;
  wire n11433_o;
  wire n11435_o;
  wire n11436_o;
  wire n11437_o;
  wire n11439_o;
  wire n11440_o;
  wire n11441_o;
  wire n11443_o;
  wire n11444_o;
  wire n11445_o;
  wire n11447_o;
  wire n11448_o;
  wire n11449_o;
  wire n11451_o;
  wire n11452_o;
  wire n11453_o;
  wire n11455_o;
  wire n11456_o;
  wire n11457_o;
  wire n11459_o;
  wire n11460_o;
  wire n11461_o;
  wire n11463_o;
  wire n11464_o;
  wire n11465_o;
  wire n11467_o;
  wire n11468_o;
  wire n11469_o;
  wire n11470_o;
  wire n11482_o;
  wire n11484_o;
  wire n11486_o;
  wire n11488_o;
  wire n11490_o;
  wire n11491_o;
  wire n11492_o;
  wire n11494_o;
  wire n11495_o;
  wire n11496_o;
  wire n11498_o;
  wire n11499_o;
  wire n11500_o;
  wire n11502_o;
  wire n11503_o;
  wire n11504_o;
  wire n11506_o;
  wire n11507_o;
  wire n11508_o;
  wire n11510_o;
  wire n11511_o;
  wire n11512_o;
  wire n11514_o;
  wire n11515_o;
  wire n11516_o;
  wire n11518_o;
  wire n11519_o;
  wire n11520_o;
  wire n11522_o;
  wire n11523_o;
  wire n11524_o;
  wire n11526_o;
  wire n11527_o;
  wire n11528_o;
  wire n11530_o;
  wire n11531_o;
  wire n11532_o;
  wire n11534_o;
  wire n11535_o;
  wire n11536_o;
  wire n11538_o;
  wire n11539_o;
  wire n11540_o;
  wire n11542_o;
  wire n11543_o;
  wire n11544_o;
  wire n11546_o;
  wire n11547_o;
  wire n11548_o;
  wire n11550_o;
  wire n11551_o;
  wire n11552_o;
  wire n11554_o;
  wire n11555_o;
  wire n11556_o;
  wire n11558_o;
  wire n11559_o;
  wire n11560_o;
  wire n11562_o;
  wire n11563_o;
  wire n11564_o;
  wire n11566_o;
  wire n11567_o;
  wire n11568_o;
  wire n11570_o;
  wire n11571_o;
  wire n11572_o;
  wire n11574_o;
  wire n11575_o;
  wire n11576_o;
  wire n11578_o;
  wire n11579_o;
  wire n11580_o;
  wire n11582_o;
  wire n11583_o;
  wire n11584_o;
  wire n11586_o;
  wire n11587_o;
  wire n11588_o;
  wire n11590_o;
  wire n11591_o;
  wire n11592_o;
  wire n11594_o;
  wire n11595_o;
  wire n11596_o;
  wire n11598_o;
  wire n11599_o;
  wire n11600_o;
  wire n11602_o;
  wire n11603_o;
  wire n11604_o;
  wire n11606_o;
  wire n11607_o;
  wire n11608_o;
  wire n11610_o;
  wire n11611_o;
  wire n11612_o;
  wire n11613_o;
  wire n11625_o;
  wire n11627_o;
  wire n11629_o;
  wire n11631_o;
  wire n11633_o;
  wire n11634_o;
  wire n11635_o;
  wire n11637_o;
  wire n11638_o;
  wire n11639_o;
  wire n11641_o;
  wire n11642_o;
  wire n11643_o;
  wire n11645_o;
  wire n11646_o;
  wire n11647_o;
  wire n11649_o;
  wire n11650_o;
  wire n11651_o;
  wire n11653_o;
  wire n11654_o;
  wire n11655_o;
  wire n11657_o;
  wire n11658_o;
  wire n11659_o;
  wire n11661_o;
  wire n11662_o;
  wire n11663_o;
  wire n11665_o;
  wire n11666_o;
  wire n11667_o;
  wire n11669_o;
  wire n11670_o;
  wire n11671_o;
  wire n11673_o;
  wire n11674_o;
  wire n11675_o;
  wire n11677_o;
  wire n11678_o;
  wire n11679_o;
  wire n11681_o;
  wire n11682_o;
  wire n11683_o;
  wire n11685_o;
  wire n11686_o;
  wire n11687_o;
  wire n11689_o;
  wire n11690_o;
  wire n11691_o;
  wire n11693_o;
  wire n11694_o;
  wire n11695_o;
  wire n11697_o;
  wire n11698_o;
  wire n11699_o;
  wire n11701_o;
  wire n11702_o;
  wire n11703_o;
  wire n11705_o;
  wire n11706_o;
  wire n11707_o;
  wire n11709_o;
  wire n11710_o;
  wire n11711_o;
  wire n11713_o;
  wire n11714_o;
  wire n11715_o;
  wire n11717_o;
  wire n11718_o;
  wire n11719_o;
  wire n11721_o;
  wire n11722_o;
  wire n11723_o;
  wire n11725_o;
  wire n11726_o;
  wire n11727_o;
  wire n11729_o;
  wire n11730_o;
  wire n11731_o;
  wire n11733_o;
  wire n11734_o;
  wire n11735_o;
  wire n11737_o;
  wire n11738_o;
  wire n11739_o;
  wire n11741_o;
  wire n11742_o;
  wire n11743_o;
  wire n11745_o;
  wire n11746_o;
  wire n11747_o;
  wire n11749_o;
  wire n11750_o;
  wire n11751_o;
  wire n11753_o;
  wire n11754_o;
  wire n11755_o;
  wire n11756_o;
  wire n11768_o;
  wire n11770_o;
  wire n11772_o;
  wire n11774_o;
  wire n11776_o;
  wire n11777_o;
  wire n11778_o;
  wire n11780_o;
  wire n11781_o;
  wire n11782_o;
  wire n11784_o;
  wire n11785_o;
  wire n11786_o;
  wire n11788_o;
  wire n11789_o;
  wire n11790_o;
  wire n11792_o;
  wire n11793_o;
  wire n11794_o;
  wire n11796_o;
  wire n11797_o;
  wire n11798_o;
  wire n11800_o;
  wire n11801_o;
  wire n11802_o;
  wire n11804_o;
  wire n11805_o;
  wire n11806_o;
  wire n11808_o;
  wire n11809_o;
  wire n11810_o;
  wire n11812_o;
  wire n11813_o;
  wire n11814_o;
  wire n11816_o;
  wire n11817_o;
  wire n11818_o;
  wire n11820_o;
  wire n11821_o;
  wire n11822_o;
  wire n11824_o;
  wire n11825_o;
  wire n11826_o;
  wire n11828_o;
  wire n11829_o;
  wire n11830_o;
  wire n11832_o;
  wire n11833_o;
  wire n11834_o;
  wire n11836_o;
  wire n11837_o;
  wire n11838_o;
  wire n11840_o;
  wire n11841_o;
  wire n11842_o;
  wire n11844_o;
  wire n11845_o;
  wire n11846_o;
  wire n11848_o;
  wire n11849_o;
  wire n11850_o;
  wire n11852_o;
  wire n11853_o;
  wire n11854_o;
  wire n11856_o;
  wire n11857_o;
  wire n11858_o;
  wire n11860_o;
  wire n11861_o;
  wire n11862_o;
  wire n11864_o;
  wire n11865_o;
  wire n11866_o;
  wire n11868_o;
  wire n11869_o;
  wire n11870_o;
  wire n11872_o;
  wire n11873_o;
  wire n11874_o;
  wire n11876_o;
  wire n11877_o;
  wire n11878_o;
  wire n11880_o;
  wire n11881_o;
  wire n11882_o;
  wire n11884_o;
  wire n11885_o;
  wire n11886_o;
  wire n11888_o;
  wire n11889_o;
  wire n11890_o;
  wire n11892_o;
  wire n11893_o;
  wire n11894_o;
  wire n11896_o;
  wire n11897_o;
  wire n11898_o;
  wire n11899_o;
  wire n11911_o;
  wire n11913_o;
  wire n11915_o;
  wire n11917_o;
  wire n11919_o;
  wire n11920_o;
  wire n11921_o;
  wire n11923_o;
  wire n11924_o;
  wire n11925_o;
  wire n11927_o;
  wire n11928_o;
  wire n11929_o;
  wire n11931_o;
  wire n11932_o;
  wire n11933_o;
  wire n11935_o;
  wire n11936_o;
  wire n11937_o;
  wire n11939_o;
  wire n11940_o;
  wire n11941_o;
  wire n11943_o;
  wire n11944_o;
  wire n11945_o;
  wire n11947_o;
  wire n11948_o;
  wire n11949_o;
  wire n11951_o;
  wire n11952_o;
  wire n11953_o;
  wire n11955_o;
  wire n11956_o;
  wire n11957_o;
  wire n11959_o;
  wire n11960_o;
  wire n11961_o;
  wire n11963_o;
  wire n11964_o;
  wire n11965_o;
  wire n11967_o;
  wire n11968_o;
  wire n11969_o;
  wire n11971_o;
  wire n11972_o;
  wire n11973_o;
  wire n11975_o;
  wire n11976_o;
  wire n11977_o;
  wire n11979_o;
  wire n11980_o;
  wire n11981_o;
  wire n11983_o;
  wire n11984_o;
  wire n11985_o;
  wire n11987_o;
  wire n11988_o;
  wire n11989_o;
  wire n11991_o;
  wire n11992_o;
  wire n11993_o;
  wire n11995_o;
  wire n11996_o;
  wire n11997_o;
  wire n11999_o;
  wire n12000_o;
  wire n12001_o;
  wire n12003_o;
  wire n12004_o;
  wire n12005_o;
  wire n12007_o;
  wire n12008_o;
  wire n12009_o;
  wire n12011_o;
  wire n12012_o;
  wire n12013_o;
  wire n12015_o;
  wire n12016_o;
  wire n12017_o;
  wire n12019_o;
  wire n12020_o;
  wire n12021_o;
  wire n12023_o;
  wire n12024_o;
  wire n12025_o;
  wire n12027_o;
  wire n12028_o;
  wire n12029_o;
  wire n12031_o;
  wire n12032_o;
  wire n12033_o;
  wire n12035_o;
  wire n12036_o;
  wire n12037_o;
  wire n12039_o;
  wire n12040_o;
  wire n12041_o;
  wire n12042_o;
  wire n12054_o;
  wire n12056_o;
  wire n12058_o;
  wire n12060_o;
  wire n12062_o;
  wire n12063_o;
  wire n12064_o;
  wire n12066_o;
  wire n12067_o;
  wire n12068_o;
  wire n12070_o;
  wire n12071_o;
  wire n12072_o;
  wire n12074_o;
  wire n12075_o;
  wire n12076_o;
  wire n12078_o;
  wire n12079_o;
  wire n12080_o;
  wire n12082_o;
  wire n12083_o;
  wire n12084_o;
  wire n12086_o;
  wire n12087_o;
  wire n12088_o;
  wire n12090_o;
  wire n12091_o;
  wire n12092_o;
  wire n12094_o;
  wire n12095_o;
  wire n12096_o;
  wire n12098_o;
  wire n12099_o;
  wire n12100_o;
  wire n12102_o;
  wire n12103_o;
  wire n12104_o;
  wire n12106_o;
  wire n12107_o;
  wire n12108_o;
  wire n12110_o;
  wire n12111_o;
  wire n12112_o;
  wire n12114_o;
  wire n12115_o;
  wire n12116_o;
  wire n12118_o;
  wire n12119_o;
  wire n12120_o;
  wire n12122_o;
  wire n12123_o;
  wire n12124_o;
  wire n12126_o;
  wire n12127_o;
  wire n12128_o;
  wire n12130_o;
  wire n12131_o;
  wire n12132_o;
  wire n12134_o;
  wire n12135_o;
  wire n12136_o;
  wire n12138_o;
  wire n12139_o;
  wire n12140_o;
  wire n12142_o;
  wire n12143_o;
  wire n12144_o;
  wire n12146_o;
  wire n12147_o;
  wire n12148_o;
  wire n12150_o;
  wire n12151_o;
  wire n12152_o;
  wire n12154_o;
  wire n12155_o;
  wire n12156_o;
  wire n12158_o;
  wire n12159_o;
  wire n12160_o;
  wire n12162_o;
  wire n12163_o;
  wire n12164_o;
  wire n12166_o;
  wire n12167_o;
  wire n12168_o;
  wire n12170_o;
  wire n12171_o;
  wire n12172_o;
  wire n12174_o;
  wire n12175_o;
  wire n12176_o;
  wire n12178_o;
  wire n12179_o;
  wire n12180_o;
  wire n12182_o;
  wire n12183_o;
  wire n12184_o;
  wire n12185_o;
  wire [3:0] n12189_o;
  wire [3:0] n12190_o;
  wire [1:0] n12191_o;
  wire [9:0] n12192_o;
  wire n12193_o;
  wire n12194_o;
  wire n12195_o;
  wire n12196_o;
  wire n12197_o;
  wire n12198_o;
  wire n12199_o;
  wire n12200_o;
  wire [3:0] n12207_o;
  wire [3:0] n12208_o;
  wire [1:0] n12209_o;
  wire [9:0] n12210_o;
  wire [2:0] n12212_o;
  wire n12218_o;
  wire n12220_o;
  wire n12222_o;
  wire n12223_o;
  wire n12224_o;
  wire n12225_o;
  wire n12226_o;
  wire n12227_o;
  wire n12228_o;
  wire n12229_o;
  wire n12230_o;
  wire n12231_o;
  wire n12232_o;
  wire n12233_o;
  wire n12234_o;
  wire n12235_o;
  wire n12236_o;
  wire n12237_o;
  wire n12238_o;
  wire n12239_o;
  wire n12240_o;
  wire [1:0] n12241_o;
  wire n12242_o;
  wire n12243_o;
  wire [2:0] n12244_o;
  wire n12245_o;
  wire [3:0] n12246_o;
  wire n12247_o;
  wire n12248_o;
  wire [4:0] n12249_o;
  wire n12250_o;
  wire [5:0] n12251_o;
  wire n12253_o;
  wire n12254_o;
  wire [1:0] n12255_o;
  wire n12256_o;
  wire [2:0] n12257_o;
  wire n12258_o;
  wire [3:0] n12259_o;
  wire n12260_o;
  wire [4:0] n12261_o;
  wire n12262_o;
  wire [5:0] n12263_o;
  wire n12269_o;
  wire n12270_o;
  wire n12271_o;
  wire n12273_o;
  wire n12275_o;
  wire n12276_o;
  wire n12277_o;
  wire n12278_o;
  wire n12279_o;
  wire n12280_o;
  wire n12281_o;
  wire n12282_o;
  wire n12283_o;
  wire n12284_o;
  wire n12285_o;
  wire n12286_o;
  wire n12287_o;
  wire n12288_o;
  wire n12289_o;
  wire n12290_o;
  wire n12291_o;
  wire n12292_o;
  wire n12293_o;
  wire n12294_o;
  wire n12295_o;
  wire n12297_o;
  wire n12298_o;
  wire [1:0] n12299_o;
  wire n12300_o;
  wire [2:0] n12301_o;
  wire n12302_o;
  wire [3:0] n12303_o;
  wire n12304_o;
  wire [4:0] n12305_o;
  wire n12306_o;
  wire [5:0] n12307_o;
  wire n12313_o;
  wire n12314_o;
  wire n12315_o;
  wire n12317_o;
  wire n12319_o;
  wire n12320_o;
  wire n12321_o;
  wire n12322_o;
  wire n12323_o;
  wire n12324_o;
  wire n12325_o;
  wire n12326_o;
  wire n12327_o;
  wire n12328_o;
  wire n12329_o;
  wire n12330_o;
  wire n12331_o;
  wire n12332_o;
  wire n12333_o;
  wire n12334_o;
  wire n12335_o;
  wire n12336_o;
  wire n12337_o;
  wire n12338_o;
  wire n12339_o;
  wire n12341_o;
  wire n12342_o;
  wire [1:0] n12343_o;
  wire n12344_o;
  wire [2:0] n12345_o;
  wire n12346_o;
  wire [3:0] n12347_o;
  wire n12348_o;
  wire [4:0] n12349_o;
  wire n12350_o;
  wire [5:0] n12351_o;
  wire n12357_o;
  wire n12358_o;
  wire n12359_o;
  wire n12361_o;
  wire n12363_o;
  wire n12364_o;
  wire n12365_o;
  wire n12366_o;
  wire n12367_o;
  wire n12368_o;
  wire n12369_o;
  wire n12370_o;
  wire n12371_o;
  wire n12372_o;
  wire n12373_o;
  wire n12374_o;
  wire n12375_o;
  wire n12376_o;
  wire n12377_o;
  wire n12378_o;
  wire n12379_o;
  wire n12380_o;
  wire n12381_o;
  wire n12382_o;
  wire n12383_o;
  wire n12385_o;
  wire n12386_o;
  wire [1:0] n12387_o;
  wire n12388_o;
  wire [2:0] n12389_o;
  wire n12390_o;
  wire [3:0] n12391_o;
  wire n12392_o;
  wire [4:0] n12393_o;
  wire n12394_o;
  wire [5:0] n12395_o;
  wire n12401_o;
  wire n12402_o;
  wire n12403_o;
  wire n12405_o;
  wire n12407_o;
  wire n12408_o;
  wire n12409_o;
  wire n12410_o;
  wire n12411_o;
  wire n12412_o;
  wire n12413_o;
  wire n12414_o;
  wire n12415_o;
  wire n12416_o;
  wire n12417_o;
  wire n12418_o;
  wire n12419_o;
  wire n12420_o;
  wire n12421_o;
  wire n12422_o;
  wire n12423_o;
  wire n12424_o;
  wire n12425_o;
  wire n12426_o;
  wire n12427_o;
  wire n12429_o;
  wire n12430_o;
  wire [1:0] n12431_o;
  wire n12432_o;
  wire [2:0] n12433_o;
  wire n12434_o;
  wire [3:0] n12435_o;
  wire n12436_o;
  wire [4:0] n12437_o;
  wire n12438_o;
  wire [5:0] n12439_o;
  wire n12445_o;
  wire n12446_o;
  wire n12447_o;
  wire n12449_o;
  wire n12451_o;
  wire n12452_o;
  wire n12453_o;
  wire n12454_o;
  wire n12455_o;
  wire n12456_o;
  wire n12457_o;
  wire n12458_o;
  wire n12459_o;
  wire n12460_o;
  wire n12461_o;
  wire n12462_o;
  wire n12463_o;
  wire n12464_o;
  wire n12465_o;
  wire n12466_o;
  wire n12467_o;
  wire n12468_o;
  wire n12469_o;
  wire n12470_o;
  wire n12471_o;
  wire n12473_o;
  wire n12474_o;
  wire [1:0] n12475_o;
  wire n12476_o;
  wire [2:0] n12477_o;
  wire n12478_o;
  wire [3:0] n12479_o;
  wire n12480_o;
  wire [4:0] n12481_o;
  wire n12482_o;
  wire [5:0] n12483_o;
  wire n12489_o;
  wire n12490_o;
  wire n12491_o;
  wire n12493_o;
  wire n12495_o;
  wire n12496_o;
  wire n12497_o;
  wire n12498_o;
  wire n12499_o;
  wire n12500_o;
  wire n12501_o;
  wire n12502_o;
  wire n12503_o;
  wire n12504_o;
  wire n12505_o;
  wire n12506_o;
  wire n12507_o;
  wire n12508_o;
  wire n12509_o;
  wire n12510_o;
  wire n12511_o;
  wire n12512_o;
  wire n12513_o;
  wire n12514_o;
  wire n12515_o;
  wire n12517_o;
  wire n12518_o;
  wire [1:0] n12519_o;
  wire n12520_o;
  wire [2:0] n12521_o;
  wire n12522_o;
  wire [3:0] n12523_o;
  wire n12524_o;
  wire [4:0] n12525_o;
  wire n12526_o;
  wire [5:0] n12527_o;
  wire n12533_o;
  wire n12534_o;
  wire n12535_o;
  wire n12537_o;
  wire n12539_o;
  wire n12540_o;
  wire n12541_o;
  wire n12542_o;
  wire n12543_o;
  wire n12544_o;
  wire n12545_o;
  wire n12546_o;
  wire n12547_o;
  wire n12548_o;
  wire n12549_o;
  wire n12550_o;
  wire n12551_o;
  wire n12552_o;
  wire n12553_o;
  wire n12554_o;
  wire n12555_o;
  wire n12556_o;
  wire n12557_o;
  wire n12558_o;
  wire n12559_o;
  wire n12561_o;
  wire n12562_o;
  wire [1:0] n12563_o;
  wire n12564_o;
  wire [2:0] n12565_o;
  wire n12566_o;
  wire [3:0] n12567_o;
  wire n12568_o;
  wire [4:0] n12569_o;
  wire n12570_o;
  wire [5:0] n12571_o;
  wire n12577_o;
  wire n12578_o;
  wire n12579_o;
  wire n12581_o;
  wire n12583_o;
  wire n12584_o;
  wire n12585_o;
  wire n12586_o;
  wire n12587_o;
  wire n12588_o;
  wire n12589_o;
  wire n12590_o;
  wire n12591_o;
  wire n12592_o;
  wire n12593_o;
  wire n12594_o;
  wire n12595_o;
  wire n12596_o;
  wire n12597_o;
  wire n12598_o;
  wire n12599_o;
  wire n12600_o;
  wire n12601_o;
  wire n12602_o;
  wire n12603_o;
  wire n12605_o;
  wire n12606_o;
  wire [1:0] n12607_o;
  wire n12608_o;
  wire [2:0] n12609_o;
  wire n12610_o;
  wire [3:0] n12611_o;
  wire n12612_o;
  wire [4:0] n12613_o;
  wire n12614_o;
  wire [5:0] n12615_o;
  wire n12621_o;
  wire n12622_o;
  wire n12623_o;
  wire n12625_o;
  wire n12627_o;
  wire n12628_o;
  wire n12629_o;
  wire n12630_o;
  wire n12631_o;
  wire n12632_o;
  wire n12633_o;
  wire n12634_o;
  wire n12635_o;
  wire n12636_o;
  wire n12637_o;
  wire n12638_o;
  wire n12639_o;
  wire n12640_o;
  wire n12641_o;
  wire n12642_o;
  wire n12643_o;
  wire n12644_o;
  wire n12645_o;
  wire n12646_o;
  wire n12647_o;
  wire n12649_o;
  wire n12650_o;
  wire [1:0] n12651_o;
  wire n12652_o;
  wire [2:0] n12653_o;
  wire n12654_o;
  wire [3:0] n12655_o;
  wire n12656_o;
  wire [4:0] n12657_o;
  wire n12658_o;
  wire [5:0] n12659_o;
  wire n12665_o;
  wire n12666_o;
  wire n12667_o;
  wire n12669_o;
  wire n12671_o;
  wire n12672_o;
  wire n12673_o;
  wire n12674_o;
  wire n12675_o;
  wire n12676_o;
  wire n12677_o;
  wire n12678_o;
  wire n12679_o;
  wire n12680_o;
  wire n12681_o;
  wire n12682_o;
  wire n12683_o;
  wire n12684_o;
  wire n12685_o;
  wire n12686_o;
  wire n12687_o;
  wire n12688_o;
  wire n12689_o;
  wire n12690_o;
  wire n12691_o;
  wire [9:0] n12692_o;
  wire [9:0] n12693_o;
  reg [9:0] regfile_block_rf0;
  reg [9:0] regfile_block_rf1;
  reg [3:0] regfile_block_rf2;
  reg [3:0] regfile_block_rf3;
  reg [2:0] regfile_block_rf4;
  reg [2:0] regfile_block_rf5;
  reg [2:0] regfile_block_rf6;
  reg [2:0] regfile_block_rf7;
  reg [2:0] regfile_block_rf8;
  reg [2:0] regfile_block_rf9;
  reg [6:0] regfile_block_rf10;
  reg [6:0] regfile_block_rf11;
  wire [30:0] regfile_block_a;
  wire [11:0] regfile_block_al;
  wire [9:0] regfile_block_nrfdo;
  wire [30:0] n12706_o;
  wire n12709_o;
  wire n12712_o;
  wire n12714_o;
  wire [3:0] n12715_o;
  wire n12717_o;
  wire [3:0] n12718_o;
  wire n12720_o;
  wire [2:0] n12721_o;
  wire n12723_o;
  wire [2:0] n12724_o;
  wire n12726_o;
  wire [2:0] n12727_o;
  wire n12729_o;
  wire [2:0] n12730_o;
  wire n12732_o;
  wire [2:0] n12733_o;
  wire n12735_o;
  wire [2:0] n12736_o;
  wire n12738_o;
  wire [6:0] n12739_o;
  wire n12741_o;
  wire [6:0] n12742_o;
  wire n12744_o;
  wire [11:0] n12745_o;
  reg [9:0] n12746_o;
  reg [9:0] n12747_o;
  reg [3:0] n12748_o;
  reg [3:0] n12749_o;
  reg [2:0] n12750_o;
  reg [2:0] n12751_o;
  reg [2:0] n12752_o;
  reg [2:0] n12753_o;
  reg [2:0] n12754_o;
  reg [2:0] n12755_o;
  reg [6:0] n12756_o;
  reg [6:0] n12757_o;
  wire [31:0] n12785_o;
  wire n12787_o;
  wire [3:0] n12788_o;
  wire [3:0] n12790_o;
  localparam [11:0] n12792_o = 12'b000000000000;
  wire [11:0] n12796_o;
  wire n12800_o;
  wire n12801_o;
  wire [1:0] n12802_o;
  wire [2:0] n12804_o;
  wire [3:0] n12806_o;
  wire [4:0] n12808_o;
  wire [5:0] n12810_o;
  wire [6:0] n12812_o;
  wire [7:0] n12814_o;
  wire [8:0] n12816_o;
  wire [9:0] n12818_o;
  wire n12819_o;
  wire [10:0] n12820_o;
  wire [11:0] n12822_o;
  wire n12828_o;
  wire n12829_o;
  wire n12830_o;
  wire n12831_o;
  wire n12833_o;
  wire n12835_o;
  wire n12836_o;
  wire n12837_o;
  wire n12838_o;
  wire n12839_o;
  wire n12840_o;
  wire n12841_o;
  wire n12842_o;
  wire n12843_o;
  wire n12844_o;
  wire n12845_o;
  wire n12846_o;
  wire n12847_o;
  wire n12848_o;
  wire n12849_o;
  wire n12850_o;
  wire n12851_o;
  wire n12852_o;
  wire n12853_o;
  wire n12854_o;
  wire n12855_o;
  wire n12856_o;
  wire n12857_o;
  wire n12858_o;
  wire n12859_o;
  wire n12860_o;
  wire n12861_o;
  wire n12862_o;
  wire n12863_o;
  wire n12864_o;
  wire n12865_o;
  wire n12866_o;
  wire n12867_o;
  wire n12868_o;
  wire n12869_o;
  wire n12870_o;
  wire n12871_o;
  wire n12872_o;
  wire n12873_o;
  wire n12874_o;
  wire n12875_o;
  wire n12876_o;
  wire n12877_o;
  wire n12878_o;
  wire n12879_o;
  wire n12880_o;
  wire n12881_o;
  wire n12882_o;
  wire n12883_o;
  wire n12884_o;
  wire n12885_o;
  wire n12886_o;
  wire n12887_o;
  wire n12888_o;
  wire n12889_o;
  wire n12890_o;
  wire n12892_o;
  wire n12893_o;
  wire [1:0] n12894_o;
  wire [2:0] n12896_o;
  wire [3:0] n12898_o;
  wire [4:0] n12900_o;
  wire [5:0] n12902_o;
  wire [6:0] n12904_o;
  wire [7:0] n12906_o;
  wire [8:0] n12908_o;
  wire [9:0] n12910_o;
  wire n12911_o;
  wire [10:0] n12912_o;
  wire [11:0] n12914_o;
  wire n12920_o;
  wire n12921_o;
  wire n12922_o;
  wire n12923_o;
  wire n12925_o;
  wire n12927_o;
  wire n12928_o;
  wire n12929_o;
  wire n12930_o;
  wire n12931_o;
  wire n12932_o;
  wire n12933_o;
  wire n12934_o;
  wire n12935_o;
  wire n12936_o;
  wire n12937_o;
  wire n12938_o;
  wire n12939_o;
  wire n12940_o;
  wire n12941_o;
  wire n12942_o;
  wire n12943_o;
  wire n12944_o;
  wire n12945_o;
  wire n12946_o;
  wire n12947_o;
  wire n12948_o;
  wire n12949_o;
  wire n12950_o;
  wire n12951_o;
  wire n12952_o;
  wire n12953_o;
  wire n12954_o;
  wire n12955_o;
  wire n12956_o;
  wire n12957_o;
  wire n12958_o;
  wire n12959_o;
  wire n12960_o;
  wire n12961_o;
  wire n12962_o;
  wire n12963_o;
  wire n12964_o;
  wire n12965_o;
  wire n12966_o;
  wire n12967_o;
  wire n12968_o;
  wire n12969_o;
  wire n12970_o;
  wire n12971_o;
  wire n12972_o;
  wire n12973_o;
  wire n12974_o;
  wire n12975_o;
  wire n12976_o;
  wire n12977_o;
  wire n12978_o;
  wire n12979_o;
  wire n12980_o;
  wire n12981_o;
  wire n12982_o;
  wire n12984_o;
  wire n12985_o;
  wire [1:0] n12986_o;
  wire [2:0] n12988_o;
  wire [3:0] n12990_o;
  wire [4:0] n12992_o;
  wire [5:0] n12994_o;
  wire [6:0] n12996_o;
  wire [7:0] n12998_o;
  wire [8:0] n13000_o;
  wire [9:0] n13002_o;
  wire n13003_o;
  wire [10:0] n13004_o;
  wire [11:0] n13006_o;
  wire n13012_o;
  wire n13013_o;
  wire n13014_o;
  wire n13015_o;
  wire n13017_o;
  wire n13019_o;
  wire n13020_o;
  wire n13021_o;
  wire n13022_o;
  wire n13023_o;
  wire n13024_o;
  wire n13025_o;
  wire n13026_o;
  wire n13027_o;
  wire n13028_o;
  wire n13029_o;
  wire n13030_o;
  wire n13031_o;
  wire n13032_o;
  wire n13033_o;
  wire n13034_o;
  wire n13035_o;
  wire n13036_o;
  wire n13037_o;
  wire n13038_o;
  wire n13039_o;
  wire n13040_o;
  wire n13041_o;
  wire n13042_o;
  wire n13043_o;
  wire n13044_o;
  wire n13045_o;
  wire n13046_o;
  wire n13047_o;
  wire n13048_o;
  wire n13049_o;
  wire n13050_o;
  wire n13051_o;
  wire n13052_o;
  wire n13053_o;
  wire n13054_o;
  wire n13055_o;
  wire n13056_o;
  wire n13057_o;
  wire n13058_o;
  wire n13059_o;
  wire n13060_o;
  wire n13061_o;
  wire n13062_o;
  wire n13063_o;
  wire n13064_o;
  wire n13065_o;
  wire n13066_o;
  wire n13067_o;
  wire n13068_o;
  wire n13069_o;
  wire n13070_o;
  wire n13071_o;
  wire n13072_o;
  wire n13073_o;
  wire n13074_o;
  wire n13076_o;
  wire n13077_o;
  wire [1:0] n13078_o;
  wire [2:0] n13080_o;
  wire [3:0] n13082_o;
  wire [4:0] n13084_o;
  wire [5:0] n13086_o;
  wire [6:0] n13088_o;
  wire [7:0] n13090_o;
  wire [8:0] n13092_o;
  wire [9:0] n13094_o;
  wire n13095_o;
  wire [10:0] n13096_o;
  wire n13097_o;
  wire [11:0] n13098_o;
  wire n13104_o;
  wire n13105_o;
  wire n13106_o;
  wire n13107_o;
  wire n13109_o;
  wire n13111_o;
  wire n13112_o;
  wire n13113_o;
  wire n13114_o;
  wire n13115_o;
  wire n13116_o;
  wire n13117_o;
  wire n13118_o;
  wire n13119_o;
  wire n13120_o;
  wire n13121_o;
  wire n13122_o;
  wire n13123_o;
  wire n13124_o;
  wire n13125_o;
  wire n13126_o;
  wire n13127_o;
  wire n13128_o;
  wire n13129_o;
  wire n13130_o;
  wire n13131_o;
  wire n13132_o;
  wire n13133_o;
  wire n13134_o;
  wire n13135_o;
  wire n13136_o;
  wire n13137_o;
  wire n13138_o;
  wire n13139_o;
  wire n13140_o;
  wire n13141_o;
  wire n13142_o;
  wire n13143_o;
  wire n13144_o;
  wire n13145_o;
  wire n13146_o;
  wire n13147_o;
  wire n13148_o;
  wire n13149_o;
  wire n13150_o;
  wire n13151_o;
  wire n13152_o;
  wire n13153_o;
  wire n13154_o;
  wire n13155_o;
  wire n13156_o;
  wire n13157_o;
  wire n13158_o;
  wire n13159_o;
  wire n13160_o;
  wire n13161_o;
  wire n13162_o;
  wire n13163_o;
  wire n13164_o;
  wire n13165_o;
  wire n13166_o;
  wire n13168_o;
  wire n13169_o;
  wire [1:0] n13170_o;
  wire [2:0] n13172_o;
  wire [3:0] n13174_o;
  wire [4:0] n13176_o;
  wire [5:0] n13178_o;
  wire [6:0] n13180_o;
  wire [7:0] n13182_o;
  wire [8:0] n13184_o;
  wire [9:0] n13186_o;
  wire n13187_o;
  wire [10:0] n13188_o;
  wire n13189_o;
  wire [11:0] n13190_o;
  wire n13196_o;
  wire n13197_o;
  wire n13198_o;
  wire n13199_o;
  wire n13201_o;
  wire n13203_o;
  wire n13204_o;
  wire n13205_o;
  wire n13206_o;
  wire n13207_o;
  wire n13208_o;
  wire n13209_o;
  wire n13210_o;
  wire n13211_o;
  wire n13212_o;
  wire n13213_o;
  wire n13214_o;
  wire n13215_o;
  wire n13216_o;
  wire n13217_o;
  wire n13218_o;
  wire n13219_o;
  wire n13220_o;
  wire n13221_o;
  wire n13222_o;
  wire n13223_o;
  wire n13224_o;
  wire n13225_o;
  wire n13226_o;
  wire n13227_o;
  wire n13228_o;
  wire n13229_o;
  wire n13230_o;
  wire n13231_o;
  wire n13232_o;
  wire n13233_o;
  wire n13234_o;
  wire n13235_o;
  wire n13236_o;
  wire n13237_o;
  wire n13238_o;
  wire n13239_o;
  wire n13240_o;
  wire n13241_o;
  wire n13242_o;
  wire n13243_o;
  wire n13244_o;
  wire n13245_o;
  wire n13246_o;
  wire n13247_o;
  wire n13248_o;
  wire n13249_o;
  wire n13250_o;
  wire n13251_o;
  wire n13252_o;
  wire n13253_o;
  wire n13254_o;
  wire n13255_o;
  wire n13256_o;
  wire n13257_o;
  wire n13258_o;
  wire n13260_o;
  wire n13261_o;
  wire [1:0] n13262_o;
  wire [2:0] n13264_o;
  wire [3:0] n13266_o;
  wire [4:0] n13268_o;
  wire [5:0] n13270_o;
  wire [6:0] n13272_o;
  wire [7:0] n13274_o;
  wire [8:0] n13276_o;
  wire [9:0] n13278_o;
  wire n13279_o;
  wire [10:0] n13280_o;
  wire n13281_o;
  wire [11:0] n13282_o;
  wire n13288_o;
  wire n13289_o;
  wire n13290_o;
  wire n13291_o;
  wire n13293_o;
  wire n13295_o;
  wire n13296_o;
  wire n13297_o;
  wire n13298_o;
  wire n13299_o;
  wire n13300_o;
  wire n13301_o;
  wire n13302_o;
  wire n13303_o;
  wire n13304_o;
  wire n13305_o;
  wire n13306_o;
  wire n13307_o;
  wire n13308_o;
  wire n13309_o;
  wire n13310_o;
  wire n13311_o;
  wire n13312_o;
  wire n13313_o;
  wire n13314_o;
  wire n13315_o;
  wire n13316_o;
  wire n13317_o;
  wire n13318_o;
  wire n13319_o;
  wire n13320_o;
  wire n13321_o;
  wire n13322_o;
  wire n13323_o;
  wire n13324_o;
  wire n13325_o;
  wire n13326_o;
  wire n13327_o;
  wire n13328_o;
  wire n13329_o;
  wire n13330_o;
  wire n13331_o;
  wire n13332_o;
  wire n13333_o;
  wire n13334_o;
  wire n13335_o;
  wire n13336_o;
  wire n13337_o;
  wire n13338_o;
  wire n13339_o;
  wire n13340_o;
  wire n13341_o;
  wire n13342_o;
  wire n13343_o;
  wire n13344_o;
  wire n13345_o;
  wire n13346_o;
  wire n13347_o;
  wire n13348_o;
  wire n13349_o;
  wire n13350_o;
  wire n13352_o;
  wire n13353_o;
  wire [1:0] n13354_o;
  wire n13355_o;
  wire [2:0] n13356_o;
  wire n13357_o;
  wire [3:0] n13358_o;
  wire [4:0] n13360_o;
  wire [5:0] n13362_o;
  wire [6:0] n13364_o;
  wire [7:0] n13366_o;
  wire [8:0] n13368_o;
  wire [9:0] n13370_o;
  wire n13371_o;
  wire [10:0] n13372_o;
  wire n13373_o;
  wire [11:0] n13374_o;
  wire n13380_o;
  wire n13381_o;
  wire n13382_o;
  wire n13383_o;
  wire n13385_o;
  wire n13387_o;
  wire n13388_o;
  wire n13389_o;
  wire n13390_o;
  wire n13391_o;
  wire n13392_o;
  wire n13393_o;
  wire n13394_o;
  wire n13395_o;
  wire n13396_o;
  wire n13397_o;
  wire n13398_o;
  wire n13399_o;
  wire n13400_o;
  wire n13401_o;
  wire n13402_o;
  wire n13403_o;
  wire n13404_o;
  wire n13405_o;
  wire n13406_o;
  wire n13407_o;
  wire n13408_o;
  wire n13409_o;
  wire n13410_o;
  wire n13411_o;
  wire n13412_o;
  wire n13413_o;
  wire n13414_o;
  wire n13415_o;
  wire n13416_o;
  wire n13417_o;
  wire n13418_o;
  wire n13419_o;
  wire n13420_o;
  wire n13421_o;
  wire n13422_o;
  wire n13423_o;
  wire n13424_o;
  wire n13425_o;
  wire n13426_o;
  wire n13427_o;
  wire n13428_o;
  wire n13429_o;
  wire n13430_o;
  wire n13431_o;
  wire n13432_o;
  wire n13433_o;
  wire n13434_o;
  wire n13435_o;
  wire n13436_o;
  wire n13437_o;
  wire n13438_o;
  wire n13439_o;
  wire n13440_o;
  wire n13441_o;
  wire n13442_o;
  wire n13444_o;
  wire n13445_o;
  wire [1:0] n13446_o;
  wire n13447_o;
  wire [2:0] n13448_o;
  wire n13449_o;
  wire [3:0] n13450_o;
  wire n13451_o;
  wire [4:0] n13452_o;
  wire n13453_o;
  wire [5:0] n13454_o;
  wire n13455_o;
  wire [6:0] n13456_o;
  wire n13457_o;
  wire [7:0] n13458_o;
  wire n13459_o;
  wire [8:0] n13460_o;
  wire n13461_o;
  wire [9:0] n13462_o;
  wire [10:0] n13464_o;
  wire n13465_o;
  wire [11:0] n13466_o;
  wire n13472_o;
  wire n13473_o;
  wire n13474_o;
  wire n13475_o;
  wire n13477_o;
  wire n13479_o;
  wire n13480_o;
  wire n13481_o;
  wire n13482_o;
  wire n13483_o;
  wire n13484_o;
  wire n13485_o;
  wire n13486_o;
  wire n13487_o;
  wire n13488_o;
  wire n13489_o;
  wire n13490_o;
  wire n13491_o;
  wire n13492_o;
  wire n13493_o;
  wire n13494_o;
  wire n13495_o;
  wire n13496_o;
  wire n13497_o;
  wire n13498_o;
  wire n13499_o;
  wire n13500_o;
  wire n13501_o;
  wire n13502_o;
  wire n13503_o;
  wire n13504_o;
  wire n13505_o;
  wire n13506_o;
  wire n13507_o;
  wire n13508_o;
  wire n13509_o;
  wire n13510_o;
  wire n13511_o;
  wire n13512_o;
  wire n13513_o;
  wire n13514_o;
  wire n13515_o;
  wire n13516_o;
  wire n13517_o;
  wire n13518_o;
  wire n13519_o;
  wire n13520_o;
  wire n13521_o;
  wire n13522_o;
  wire n13523_o;
  wire n13524_o;
  wire n13525_o;
  wire n13526_o;
  wire n13527_o;
  wire n13528_o;
  wire n13529_o;
  wire n13530_o;
  wire n13531_o;
  wire n13532_o;
  wire n13533_o;
  wire n13534_o;
  wire n13536_o;
  wire n13537_o;
  wire [1:0] n13538_o;
  wire n13539_o;
  wire [2:0] n13540_o;
  wire n13541_o;
  wire [3:0] n13542_o;
  wire n13543_o;
  wire [4:0] n13544_o;
  wire n13545_o;
  wire [5:0] n13546_o;
  wire n13547_o;
  wire [6:0] n13548_o;
  wire n13549_o;
  wire [7:0] n13550_o;
  wire n13551_o;
  wire [8:0] n13552_o;
  wire n13553_o;
  wire [9:0] n13554_o;
  wire [10:0] n13556_o;
  wire n13557_o;
  wire [11:0] n13558_o;
  wire n13564_o;
  wire n13565_o;
  wire n13566_o;
  wire n13567_o;
  wire n13569_o;
  wire n13571_o;
  wire n13572_o;
  wire n13573_o;
  wire n13574_o;
  wire n13575_o;
  wire n13576_o;
  wire n13577_o;
  wire n13578_o;
  wire n13579_o;
  wire n13580_o;
  wire n13581_o;
  wire n13582_o;
  wire n13583_o;
  wire n13584_o;
  wire n13585_o;
  wire n13586_o;
  wire n13587_o;
  wire n13588_o;
  wire n13589_o;
  wire n13590_o;
  wire n13591_o;
  wire n13592_o;
  wire n13593_o;
  wire n13594_o;
  wire n13595_o;
  wire n13596_o;
  wire n13597_o;
  wire n13598_o;
  wire n13599_o;
  wire n13600_o;
  wire n13601_o;
  wire n13602_o;
  wire n13603_o;
  wire n13604_o;
  wire n13605_o;
  wire n13606_o;
  wire n13607_o;
  wire n13608_o;
  wire n13609_o;
  wire n13610_o;
  wire n13611_o;
  wire n13612_o;
  wire n13613_o;
  wire n13614_o;
  wire n13615_o;
  wire n13616_o;
  wire n13617_o;
  wire n13618_o;
  wire n13619_o;
  wire n13620_o;
  wire n13621_o;
  wire n13622_o;
  wire n13623_o;
  wire n13624_o;
  wire n13625_o;
  wire n13626_o;
  wire n13628_o;
  wire n13629_o;
  wire [1:0] n13630_o;
  wire n13631_o;
  wire [2:0] n13632_o;
  wire n13633_o;
  wire [3:0] n13634_o;
  wire n13635_o;
  wire [4:0] n13636_o;
  wire n13637_o;
  wire [5:0] n13638_o;
  wire n13639_o;
  wire [6:0] n13640_o;
  wire n13641_o;
  wire [7:0] n13642_o;
  wire n13643_o;
  wire [8:0] n13644_o;
  wire n13645_o;
  wire [9:0] n13646_o;
  wire [10:0] n13648_o;
  wire n13649_o;
  wire [11:0] n13650_o;
  wire n13656_o;
  wire n13657_o;
  wire n13658_o;
  wire n13659_o;
  wire n13661_o;
  wire n13663_o;
  wire n13664_o;
  wire n13665_o;
  wire n13666_o;
  wire n13667_o;
  wire n13668_o;
  wire n13669_o;
  wire n13670_o;
  wire n13671_o;
  wire n13672_o;
  wire n13673_o;
  wire n13674_o;
  wire n13675_o;
  wire n13676_o;
  wire n13677_o;
  wire n13678_o;
  wire n13679_o;
  wire n13680_o;
  wire n13681_o;
  wire n13682_o;
  wire n13683_o;
  wire n13684_o;
  wire n13685_o;
  wire n13686_o;
  wire n13687_o;
  wire n13688_o;
  wire n13689_o;
  wire n13690_o;
  wire n13691_o;
  wire n13692_o;
  wire n13693_o;
  wire n13694_o;
  wire n13695_o;
  wire n13696_o;
  wire n13697_o;
  wire n13698_o;
  wire n13699_o;
  wire n13700_o;
  wire n13701_o;
  wire n13702_o;
  wire n13703_o;
  wire n13704_o;
  wire n13705_o;
  wire n13706_o;
  wire n13707_o;
  wire n13708_o;
  wire n13709_o;
  wire n13710_o;
  wire n13711_o;
  wire n13712_o;
  wire n13713_o;
  wire n13714_o;
  wire n13715_o;
  wire n13716_o;
  wire n13717_o;
  wire n13718_o;
  wire [9:0] n13719_o;
  wire [2:0] n13721_o;
  wire n13727_o;
  wire n13729_o;
  wire n13731_o;
  wire n13732_o;
  wire n13733_o;
  wire n13734_o;
  wire n13735_o;
  wire [9:0] n13736_o;
  reg [9:0] n13737_q;
  wire [9:0] n13738_o;
  reg [9:0] n13739_q;
  wire [3:0] n13740_o;
  reg [3:0] n13741_q;
  wire [3:0] n13742_o;
  reg [3:0] n13743_q;
  wire [2:0] n13744_o;
  reg [2:0] n13745_q;
  wire [2:0] n13746_o;
  reg [2:0] n13747_q;
  wire [2:0] n13748_o;
  reg [2:0] n13749_q;
  wire [2:0] n13750_o;
  reg [2:0] n13751_q;
  wire [2:0] n13752_o;
  reg [2:0] n13753_q;
  wire [2:0] n13754_o;
  reg [2:0] n13755_q;
  wire [6:0] n13756_o;
  reg [6:0] n13757_q;
  wire [6:0] n13758_o;
  reg [6:0] n13759_q;
  wire [9:0] n13760_o;
  wire [9:0] addshift_block_nidlat;
  wire [9:0] addshift_block_port_nid;
  wire [9:0] addshift_block_port_rf;
  wire [11:0] addshift_block_sumlat;
  wire [10:0] addshift_block_cin;
  wire [10:0] addshift_block_sum;
  wire addshift_block_idpos;
  wire n13762_o;
  wire n13763_o;
  wire n13768_o;
  wire n13769_o;
  wire n13770_o;
  wire n13771_o;
  wire n13774_o;
  wire n13781_o;
  wire n13782_o;
  wire n13788_o;
  wire n13789_o;
  wire n13790_o;
  wire n13791_o;
  wire n13792_o;
  wire n13798_o;
  wire n13799_o;
  wire n13800_o;
  wire n13801_o;
  wire n13802_o;
  wire n13803_o;
  wire n13804_o;
  wire n13805_o;
  wire n13806_o;
  wire n13807_o;
  wire n13808_o;
  wire n13809_o;
  wire n13810_o;
  wire n13811_o;
  wire n13812_o;
  wire n13813_o;
  wire n13814_o;
  wire n13815_o;
  wire n13816_o;
  wire n13817_o;
  wire n13818_o;
  wire n13821_o;
  wire n13828_o;
  wire n13829_o;
  wire n13837_o;
  wire n13844_o;
  wire n13845_o;
  wire n13851_o;
  wire n13852_o;
  wire n13853_o;
  wire n13854_o;
  wire n13855_o;
  wire n13861_o;
  wire n13862_o;
  wire n13863_o;
  wire n13864_o;
  wire n13865_o;
  wire n13866_o;
  wire n13867_o;
  wire n13868_o;
  wire n13869_o;
  wire n13870_o;
  wire n13871_o;
  wire n13872_o;
  wire n13873_o;
  wire n13874_o;
  wire n13875_o;
  wire n13876_o;
  wire n13877_o;
  wire n13878_o;
  wire n13879_o;
  wire n13880_o;
  wire n13881_o;
  wire n13884_o;
  wire n13891_o;
  wire n13892_o;
  wire n13900_o;
  wire n13907_o;
  wire n13908_o;
  wire n13914_o;
  wire n13915_o;
  wire n13916_o;
  wire n13917_o;
  wire n13918_o;
  wire n13924_o;
  wire n13925_o;
  wire n13926_o;
  wire n13927_o;
  wire n13928_o;
  wire n13929_o;
  wire n13930_o;
  wire n13931_o;
  wire n13932_o;
  wire n13933_o;
  wire n13934_o;
  wire n13935_o;
  wire n13936_o;
  wire n13937_o;
  wire n13938_o;
  wire n13939_o;
  wire n13940_o;
  wire n13941_o;
  wire n13942_o;
  wire n13943_o;
  wire n13944_o;
  wire n13947_o;
  wire n13954_o;
  wire n13955_o;
  wire n13963_o;
  wire n13970_o;
  wire n13971_o;
  wire n13977_o;
  wire n13978_o;
  wire n13979_o;
  wire n13980_o;
  wire n13981_o;
  wire n13987_o;
  wire n13988_o;
  wire n13989_o;
  wire n13990_o;
  wire n13991_o;
  wire n13992_o;
  wire n13993_o;
  wire n13994_o;
  wire n13995_o;
  wire n13996_o;
  wire n13997_o;
  wire n13998_o;
  wire n13999_o;
  wire n14000_o;
  wire n14001_o;
  wire n14002_o;
  wire n14003_o;
  wire n14004_o;
  wire n14005_o;
  wire n14006_o;
  wire n14007_o;
  wire n14010_o;
  wire n14017_o;
  wire n14018_o;
  wire n14026_o;
  wire n14033_o;
  wire n14034_o;
  wire n14040_o;
  wire n14041_o;
  wire n14042_o;
  wire n14043_o;
  wire n14044_o;
  wire n14050_o;
  wire n14051_o;
  wire n14052_o;
  wire n14053_o;
  wire n14054_o;
  wire n14055_o;
  wire n14056_o;
  wire n14057_o;
  wire n14058_o;
  wire n14059_o;
  wire n14060_o;
  wire n14061_o;
  wire n14062_o;
  wire n14063_o;
  wire n14064_o;
  wire n14065_o;
  wire n14066_o;
  wire n14067_o;
  wire n14068_o;
  wire n14069_o;
  wire n14070_o;
  wire n14073_o;
  wire n14080_o;
  wire n14081_o;
  wire n14089_o;
  wire n14096_o;
  wire n14097_o;
  wire n14103_o;
  wire n14104_o;
  wire n14105_o;
  wire n14106_o;
  wire n14107_o;
  wire n14113_o;
  wire n14114_o;
  wire n14115_o;
  wire n14116_o;
  wire n14117_o;
  wire n14118_o;
  wire n14119_o;
  wire n14120_o;
  wire n14121_o;
  wire n14122_o;
  wire n14123_o;
  wire n14124_o;
  wire n14125_o;
  wire n14126_o;
  wire n14127_o;
  wire n14128_o;
  wire n14129_o;
  wire n14130_o;
  wire n14131_o;
  wire n14132_o;
  wire n14133_o;
  wire n14136_o;
  wire n14143_o;
  wire n14144_o;
  wire n14152_o;
  wire n14159_o;
  wire n14160_o;
  wire n14166_o;
  wire n14167_o;
  wire n14168_o;
  wire n14169_o;
  wire n14170_o;
  wire n14176_o;
  wire n14177_o;
  wire n14178_o;
  wire n14179_o;
  wire n14180_o;
  wire n14181_o;
  wire n14182_o;
  wire n14183_o;
  wire n14184_o;
  wire n14185_o;
  wire n14186_o;
  wire n14187_o;
  wire n14188_o;
  wire n14189_o;
  wire n14190_o;
  wire n14191_o;
  wire n14192_o;
  wire n14193_o;
  wire n14194_o;
  wire n14195_o;
  wire n14196_o;
  wire n14199_o;
  wire n14206_o;
  wire n14207_o;
  wire n14215_o;
  wire n14222_o;
  wire n14223_o;
  wire n14229_o;
  wire n14230_o;
  wire n14231_o;
  wire n14232_o;
  wire n14233_o;
  wire n14239_o;
  wire n14240_o;
  wire n14241_o;
  wire n14242_o;
  wire n14243_o;
  wire n14244_o;
  wire n14245_o;
  wire n14246_o;
  wire n14247_o;
  wire n14248_o;
  wire n14249_o;
  wire n14250_o;
  wire n14251_o;
  wire n14252_o;
  wire n14253_o;
  wire n14254_o;
  wire n14255_o;
  wire n14256_o;
  wire n14257_o;
  wire n14258_o;
  wire n14259_o;
  wire n14262_o;
  wire n14269_o;
  wire n14270_o;
  wire n14278_o;
  wire n14285_o;
  wire n14286_o;
  wire n14292_o;
  wire n14293_o;
  wire n14294_o;
  wire n14295_o;
  wire n14296_o;
  wire n14302_o;
  wire n14303_o;
  wire n14304_o;
  wire n14305_o;
  wire n14306_o;
  wire n14307_o;
  wire n14308_o;
  wire n14309_o;
  wire n14310_o;
  wire n14311_o;
  wire n14312_o;
  wire n14313_o;
  wire n14314_o;
  wire n14315_o;
  wire n14316_o;
  wire n14317_o;
  wire n14318_o;
  wire n14319_o;
  wire n14320_o;
  wire n14321_o;
  wire n14322_o;
  wire n14325_o;
  wire n14332_o;
  wire n14333_o;
  wire n14341_o;
  wire n14348_o;
  wire n14349_o;
  wire n14355_o;
  wire n14356_o;
  wire n14357_o;
  wire n14358_o;
  wire n14359_o;
  wire n14365_o;
  wire n14366_o;
  wire n14367_o;
  wire n14368_o;
  wire n14369_o;
  wire n14370_o;
  wire n14371_o;
  wire n14372_o;
  wire n14373_o;
  wire n14374_o;
  wire n14375_o;
  wire n14376_o;
  wire n14377_o;
  wire n14378_o;
  wire n14379_o;
  wire n14380_o;
  wire n14381_o;
  wire n14382_o;
  wire n14383_o;
  wire n14384_o;
  wire n14385_o;
  wire n14388_o;
  wire n14395_o;
  wire n14396_o;
  wire n14402_o;
  wire n14403_o;
  wire n14404_o;
  wire n14405_o;
  wire n14406_o;
  wire n14409_o;
  wire n14416_o;
  wire n14417_o;
  wire n14423_o;
  wire [9:0] n14424_o;
  wire n14425_o;
  wire n14426_o;
  reg n14427_q;
  wire n14428_o;
  wire n14429_o;
  reg n14430_q;
  wire n14431_o;
  wire n14432_o;
  reg n14433_q;
  wire n14434_o;
  wire n14435_o;
  reg n14436_q;
  wire n14437_o;
  wire n14438_o;
  reg n14439_q;
  wire n14440_o;
  wire n14441_o;
  reg n14442_q;
  wire n14443_o;
  wire n14444_o;
  reg n14445_q;
  wire n14446_o;
  wire n14447_o;
  reg n14448_q;
  wire n14449_o;
  wire n14450_o;
  reg n14451_q;
  wire n14452_o;
  wire n14453_o;
  reg n14454_q;
  wire [9:0] n14455_o;
  wire [9:0] n14456_o;
  wire [9:0] n14457_o;
  wire n14458_o;
  wire n14459_o;
  reg n14460_q;
  wire n14461_o;
  wire n14462_o;
  reg n14463_q;
  wire n14464_o;
  wire n14465_o;
  reg n14466_q;
  wire n14467_o;
  wire n14468_o;
  reg n14469_q;
  wire n14470_o;
  wire n14471_o;
  reg n14472_q;
  wire n14473_o;
  wire n14474_o;
  reg n14475_q;
  wire n14476_o;
  wire n14477_o;
  reg n14478_q;
  wire n14479_o;
  wire n14480_o;
  reg n14481_q;
  wire n14482_o;
  wire n14483_o;
  reg n14484_q;
  wire n14485_o;
  wire n14486_o;
  reg n14487_q;
  wire n14488_o;
  wire n14489_o;
  reg n14490_q;
  wire [11:0] n14491_o;
  wire [10:0] n14492_o;
  wire [10:0] n14493_o;
  reg [6:0] pitchinc_block_pitchlat;
  reg [6:0] pitchinc_block_pitchreg;
  wire [7:0] pitchinc_block_toggle;
  wire n14502_o;
  wire n14503_o;
  wire n14504_o;
  wire n14505_o;
  wire n14506_o;
  wire n14507_o;
  wire n14508_o;
  wire [3:0] n14509_o;
  wire n14514_o;
  wire n14515_o;
  wire n14516_o;
  wire n14517_o;
  wire n14518_o;
  wire [3:0] n14519_o;
  wire n14522_o;
  wire n14529_o;
  wire [6:0] n14530_o;
  wire n14541_o;
  wire n14543_o;
  wire n14545_o;
  wire n14546_o;
  wire n14547_o;
  wire n14548_o;
  wire n14549_o;
  wire n14550_o;
  wire n14551_o;
  wire n14552_o;
  wire n14553_o;
  wire n14554_o;
  wire n14555_o;
  wire n14556_o;
  wire n14557_o;
  wire n14558_o;
  wire n14559_o;
  wire n14560_o;
  wire n14561_o;
  wire n14562_o;
  wire n14563_o;
  wire n14564_o;
  wire n14565_o;
  wire n14566_o;
  wire n14567_o;
  wire n14568_o;
  wire n14569_o;
  wire n14570_o;
  wire n14571_o;
  wire n14572_o;
  wire n14573_o;
  wire n14574_o;
  wire n14575_o;
  wire n14576_o;
  wire n14577_o;
  wire n14578_o;
  wire n14579_o;
  wire [6:0] n14580_o;
  wire [6:0] n14581_o;
  wire n14587_o;
  wire n14588_o;
  wire n14589_o;
  wire n14590_o;
  wire n14591_o;
  wire n14592_o;
  wire n14593_o;
  wire n14594_o;
  wire n14595_o;
  wire n14596_o;
  wire n14597_o;
  wire n14598_o;
  wire n14599_o;
  wire n14600_o;
  wire n14601_o;
  wire n14602_o;
  wire n14603_o;
  wire n14604_o;
  wire n14605_o;
  wire n14606_o;
  wire n14607_o;
  wire n14608_o;
  wire n14609_o;
  wire n14610_o;
  wire n14611_o;
  wire n14612_o;
  wire n14613_o;
  wire n14614_o;
  wire n14615_o;
  wire n14616_o;
  wire n14617_o;
  wire n14618_o;
  wire n14619_o;
  wire n14620_o;
  wire n14621_o;
  wire n14622_o;
  wire [6:0] n14623_o;
  reg [6:0] n14624_q;
  wire [6:0] n14625_o;
  reg [6:0] n14626_q;
  wire [7:0] n14627_o;
  wire n14629_o;
  wire n14630_o;
  wire n14631_o;
  wire n14632_o;
  wire n14633_o;
  wire n14638_o;
  wire n14639_o;
  wire n14640_o;
  wire [5:0] nid_block_wl;
  wire [1:0] n14641_o;
  wire [2:0] n14642_o;
  wire [3:0] n14643_o;
  wire [4:0] n14644_o;
  wire [5:0] n14645_o;
  wire n14647_o;
  wire n14648_o;
  wire [1:0] n14649_o;
  wire n14650_o;
  wire [2:0] n14651_o;
  wire [3:0] n14653_o;
  wire n14654_o;
  wire n14655_o;
  wire [4:0] n14656_o;
  wire n14657_o;
  wire [5:0] n14658_o;
  wire n14664_o;
  wire n14665_o;
  wire n14666_o;
  wire n14668_o;
  wire n14670_o;
  wire n14671_o;
  wire n14672_o;
  wire n14673_o;
  wire n14674_o;
  wire n14675_o;
  wire n14676_o;
  wire n14677_o;
  wire n14678_o;
  wire n14679_o;
  wire n14680_o;
  wire n14681_o;
  wire n14682_o;
  wire n14683_o;
  wire n14684_o;
  wire n14685_o;
  wire n14686_o;
  wire n14687_o;
  wire n14688_o;
  wire n14689_o;
  wire n14690_o;
  wire n14692_o;
  wire n14693_o;
  wire [1:0] n14694_o;
  wire n14695_o;
  wire [2:0] n14696_o;
  wire [3:0] n14698_o;
  wire n14699_o;
  wire n14700_o;
  wire [4:0] n14701_o;
  wire n14702_o;
  wire [5:0] n14703_o;
  wire n14709_o;
  wire n14710_o;
  wire n14711_o;
  wire n14713_o;
  wire n14715_o;
  wire n14716_o;
  wire n14717_o;
  wire n14718_o;
  wire n14719_o;
  wire n14720_o;
  wire n14721_o;
  wire n14722_o;
  wire n14723_o;
  wire n14724_o;
  wire n14725_o;
  wire n14726_o;
  wire n14727_o;
  wire n14728_o;
  wire n14729_o;
  wire n14730_o;
  wire n14731_o;
  wire n14732_o;
  wire n14733_o;
  wire n14734_o;
  wire n14735_o;
  wire n14737_o;
  wire n14738_o;
  wire [1:0] n14739_o;
  wire n14740_o;
  wire [2:0] n14741_o;
  wire [3:0] n14743_o;
  wire n14744_o;
  wire n14745_o;
  wire [4:0] n14746_o;
  wire n14747_o;
  wire [5:0] n14748_o;
  wire n14754_o;
  wire n14755_o;
  wire n14756_o;
  wire n14758_o;
  wire n14760_o;
  wire n14761_o;
  wire n14762_o;
  wire n14763_o;
  wire n14764_o;
  wire n14765_o;
  wire n14766_o;
  wire n14767_o;
  wire n14768_o;
  wire n14769_o;
  wire n14770_o;
  wire n14771_o;
  wire n14772_o;
  wire n14773_o;
  wire n14774_o;
  wire n14775_o;
  wire n14776_o;
  wire n14777_o;
  wire n14778_o;
  wire n14779_o;
  wire n14780_o;
  wire n14782_o;
  wire n14783_o;
  wire [1:0] n14784_o;
  wire n14785_o;
  wire [2:0] n14786_o;
  wire [3:0] n14788_o;
  wire n14789_o;
  wire n14790_o;
  wire [4:0] n14791_o;
  wire n14792_o;
  wire [5:0] n14793_o;
  wire n14799_o;
  wire n14800_o;
  wire n14801_o;
  wire n14803_o;
  wire n14805_o;
  wire n14806_o;
  wire n14807_o;
  wire n14808_o;
  wire n14809_o;
  wire n14810_o;
  wire n14811_o;
  wire n14812_o;
  wire n14813_o;
  wire n14814_o;
  wire n14815_o;
  wire n14816_o;
  wire n14817_o;
  wire n14818_o;
  wire n14819_o;
  wire n14820_o;
  wire n14821_o;
  wire n14822_o;
  wire n14823_o;
  wire n14824_o;
  wire n14825_o;
  wire n14827_o;
  wire n14828_o;
  wire [1:0] n14829_o;
  wire n14830_o;
  wire [2:0] n14831_o;
  wire [3:0] n14833_o;
  wire n14834_o;
  wire n14835_o;
  wire [4:0] n14836_o;
  wire n14837_o;
  wire [5:0] n14838_o;
  wire n14844_o;
  wire n14845_o;
  wire n14846_o;
  wire n14848_o;
  wire n14850_o;
  wire n14851_o;
  wire n14852_o;
  wire n14853_o;
  wire n14854_o;
  wire n14855_o;
  wire n14856_o;
  wire n14857_o;
  wire n14858_o;
  wire n14859_o;
  wire n14860_o;
  wire n14861_o;
  wire n14862_o;
  wire n14863_o;
  wire n14864_o;
  wire n14865_o;
  wire n14866_o;
  wire n14867_o;
  wire n14868_o;
  wire n14869_o;
  wire n14870_o;
  wire n14872_o;
  wire n14873_o;
  wire [1:0] n14874_o;
  wire n14875_o;
  wire [2:0] n14876_o;
  wire [3:0] n14878_o;
  wire n14879_o;
  wire n14880_o;
  wire [4:0] n14881_o;
  wire n14882_o;
  wire [5:0] n14883_o;
  wire n14889_o;
  wire n14890_o;
  wire n14891_o;
  wire n14893_o;
  wire n14895_o;
  wire n14896_o;
  wire n14897_o;
  wire n14898_o;
  wire n14899_o;
  wire n14900_o;
  wire n14901_o;
  wire n14902_o;
  wire n14903_o;
  wire n14904_o;
  wire n14905_o;
  wire n14906_o;
  wire n14907_o;
  wire n14908_o;
  wire n14909_o;
  wire n14910_o;
  wire n14911_o;
  wire n14912_o;
  wire n14913_o;
  wire n14914_o;
  wire n14915_o;
  wire n14917_o;
  wire n14918_o;
  wire [1:0] n14919_o;
  wire n14920_o;
  wire [2:0] n14921_o;
  wire [3:0] n14922_o;
  wire n14923_o;
  wire n14924_o;
  wire [4:0] n14925_o;
  wire n14926_o;
  wire [5:0] n14927_o;
  wire n14933_o;
  wire n14934_o;
  wire n14935_o;
  wire n14937_o;
  wire n14939_o;
  wire n14940_o;
  wire n14941_o;
  wire n14942_o;
  wire n14943_o;
  wire n14944_o;
  wire n14945_o;
  wire n14946_o;
  wire n14947_o;
  wire n14948_o;
  wire n14949_o;
  wire n14950_o;
  wire n14951_o;
  wire n14952_o;
  wire n14953_o;
  wire n14954_o;
  wire n14955_o;
  wire n14956_o;
  wire n14957_o;
  wire n14958_o;
  wire n14959_o;
  wire n14961_o;
  wire n14962_o;
  wire [1:0] n14963_o;
  wire n14964_o;
  wire [2:0] n14965_o;
  wire [3:0] n14967_o;
  wire n14968_o;
  wire n14969_o;
  wire [4:0] n14970_o;
  wire n14971_o;
  wire [5:0] n14972_o;
  wire n14978_o;
  wire n14979_o;
  wire n14980_o;
  wire n14982_o;
  wire n14984_o;
  wire n14985_o;
  wire n14986_o;
  wire n14987_o;
  wire n14988_o;
  wire n14989_o;
  wire n14990_o;
  wire n14991_o;
  wire n14992_o;
  wire n14993_o;
  wire n14994_o;
  wire n14995_o;
  wire n14996_o;
  wire n14997_o;
  wire n14998_o;
  wire n14999_o;
  wire n15000_o;
  wire n15001_o;
  wire n15002_o;
  wire n15003_o;
  wire n15004_o;
  wire n15006_o;
  wire n15007_o;
  wire [1:0] n15008_o;
  wire n15009_o;
  wire [2:0] n15010_o;
  wire [3:0] n15012_o;
  wire [4:0] n15014_o;
  wire n15015_o;
  wire [5:0] n15016_o;
  wire n15022_o;
  wire n15023_o;
  wire n15024_o;
  wire n15026_o;
  wire n15028_o;
  wire n15029_o;
  wire n15030_o;
  wire n15031_o;
  wire n15032_o;
  wire n15033_o;
  wire n15034_o;
  wire n15035_o;
  wire n15036_o;
  wire n15037_o;
  wire n15038_o;
  wire n15039_o;
  wire n15040_o;
  wire n15041_o;
  wire n15042_o;
  wire n15043_o;
  wire n15044_o;
  wire n15045_o;
  wire n15046_o;
  wire n15047_o;
  wire n15048_o;
  wire n15050_o;
  wire n15051_o;
  wire [1:0] n15052_o;
  wire n15053_o;
  wire [2:0] n15054_o;
  wire [3:0] n15056_o;
  wire [4:0] n15058_o;
  wire n15059_o;
  wire [5:0] n15060_o;
  wire n15066_o;
  wire n15067_o;
  wire n15068_o;
  wire n15070_o;
  wire n15072_o;
  wire n15073_o;
  wire n15074_o;
  wire n15075_o;
  wire n15076_o;
  wire n15077_o;
  wire n15078_o;
  wire n15079_o;
  wire n15080_o;
  wire n15081_o;
  wire n15082_o;
  wire n15083_o;
  wire n15084_o;
  wire n15085_o;
  wire n15086_o;
  wire n15087_o;
  wire n15088_o;
  wire n15089_o;
  wire n15090_o;
  wire n15091_o;
  wire n15092_o;
  wire idlat_block_idlaten;
  wire idlat_block_n;
  wire n15094_o;
  wire n15095_o;
  wire n15096_o;
  wire n15097_o;
  wire n15098_o;
  wire n15103_o;
  wire n15104_o;
  wire n15105_o;
  wire n15107_o;
  wire n15108_o;
  wire n15109_o;
  wire n15114_o;
  wire n15115_o;
  wire n15116_o;
  wire n15118_o;
  wire n15123_o;
  wire n15124_o;
  wire n15125_o;
  wire n15126_o;
  wire n15127_o;
  wire n15128_o;
  wire n15129_o;
  wire n15130_o;
  wire n15131_o;
  wire n15132_o;
  wire n15133_o;
  wire n15134_o;
  wire n15135_o;
  wire n15138_o;
  wire [7:0] n15140_o;
  wire [7:0] n15145_o;
  wire n15151_o;
  wire n15153_o;
  wire n15155_o;
  wire n15156_o;
  wire n15157_o;
  wire n15158_o;
  wire n15159_o;
  wire n15160_o;
  wire n15161_o;
  wire n15162_o;
  wire n15163_o;
  wire n15164_o;
  wire n15165_o;
  wire n15166_o;
  wire n15167_o;
  wire n15168_o;
  wire n15169_o;
  wire [3:0] mem_block_swapa;
  wire [30:0] mem_block_a;
  wire mem_block_clkmem0;
  wire mem_block_clkmem1;
  wire mem_block_clkmem2;
  wire n15173_o;
  wire n15174_o;
  wire n15175_o;
  wire n15176_o;
  wire [30:0] n15177_o;
  wire n15179_o;
  wire n15180_o;
  wire n15181_o;
  wire n15182_o;
  wire n15183_o;
  wire n15184_o;
  wire n15185_o;
  wire n15190_o;
  wire n15191_o;
  wire n15192_o;
  wire n15194_o;
  wire n15195_o;
  wire n15196_o;
  wire n15201_o;
  wire n15202_o;
  wire n15203_o;
  wire n15205_o;
  wire [31:0] n15207_o;
  wire n15209_o;
  wire [3:0] n15210_o;
  wire n15216_o;
  wire [3:0] n15219_o;
  wire [9:0] n15224_o;
  wire [31:0] n15225_o;
  wire n15227_o;
  wire [9:0] n15228_o;
  wire [9:0] n15230_o;
  wire n15232_o;
  wire n15237_o;
  wire n15238_o;
  wire n15240_o;
  wire n15241_o;
  wire n15246_o;
  wire n15247_o;
  wire n15248_o;
  wire n15250_o;
  wire [31:0] n15252_o;
  wire n15254_o;
  wire [3:0] n15255_o;
  wire n15261_o;
  wire [3:0] n15264_o;
  wire [11:0] n15269_o;
  wire [31:0] n15270_o;
  wire n15272_o;
  wire [11:0] n15273_o;
  wire n15276_o;
  wire n15281_o;
  wire n15282_o;
  wire n15284_o;
  wire n15285_o;
  wire n15286_o;
  wire n15291_o;
  wire n15292_o;
  wire n15293_o;
  wire n15295_o;
  wire [31:0] n15297_o;
  wire n15299_o;
  wire [3:0] n15300_o;
  wire n15306_o;
  wire [3:0] n15309_o;
  wire [11:0] n15314_o;
  wire [31:0] n15315_o;
  wire n15317_o;
  wire [11:0] n15318_o;
  wire [3:0] n15320_o;
  wire [11:0] arithmetic_block_memxdo;
  wire [1:0] arithmetic_block_wl;
  wire [57:0] arithmetic_block_row0;
  wire [57:0] arithmetic_block_row1;
  wire [57:0] arithmetic_block_row2;
  wire [57:0] arithmetic_block_row3;
  wire [57:0] arithmetic_block_row4;
  wire [11:0] arithmetic_block_memlatmuxq;
  wire [23:0] arithmetic_block_memlatmux;
  wire [48:0] arithmetic_block_iereg;
  wire n15327_o;
  wire n15328_o;
  wire n15329_o;
  wire [1:0] n15330_o;
  wire n15332_o;
  wire n15333_o;
  wire [1:0] n15334_o;
  wire n15340_o;
  wire n15341_o;
  wire n15342_o;
  wire n15344_o;
  wire n15346_o;
  wire n15347_o;
  wire n15348_o;
  wire n15349_o;
  wire n15350_o;
  wire n15352_o;
  wire n15353_o;
  wire [1:0] n15354_o;
  wire n15360_o;
  wire n15361_o;
  wire n15362_o;
  wire n15364_o;
  wire n15366_o;
  wire n15367_o;
  wire n15368_o;
  wire n15369_o;
  wire n15370_o;
  wire n15372_o;
  wire n15373_o;
  wire [1:0] n15374_o;
  wire n15380_o;
  wire n15381_o;
  wire n15382_o;
  wire n15384_o;
  wire n15386_o;
  wire n15387_o;
  wire n15388_o;
  wire n15389_o;
  wire n15390_o;
  wire n15392_o;
  wire n15393_o;
  wire [1:0] n15394_o;
  wire n15400_o;
  wire n15401_o;
  wire n15402_o;
  wire n15404_o;
  wire n15406_o;
  wire n15407_o;
  wire n15408_o;
  wire n15409_o;
  wire n15410_o;
  wire n15412_o;
  wire n15413_o;
  wire [1:0] n15414_o;
  wire n15420_o;
  wire n15421_o;
  wire n15422_o;
  wire n15424_o;
  wire n15426_o;
  wire n15427_o;
  wire n15428_o;
  wire n15429_o;
  wire n15430_o;
  wire n15432_o;
  wire n15433_o;
  wire [1:0] n15434_o;
  wire n15440_o;
  wire n15441_o;
  wire n15442_o;
  wire n15444_o;
  wire n15446_o;
  wire n15447_o;
  wire n15448_o;
  wire n15449_o;
  wire n15450_o;
  wire n15452_o;
  wire n15453_o;
  wire [1:0] n15454_o;
  wire n15460_o;
  wire n15461_o;
  wire n15462_o;
  wire n15464_o;
  wire n15466_o;
  wire n15467_o;
  wire n15468_o;
  wire n15469_o;
  wire n15470_o;
  wire n15472_o;
  wire n15473_o;
  wire [1:0] n15474_o;
  wire n15480_o;
  wire n15481_o;
  wire n15482_o;
  wire n15484_o;
  wire n15486_o;
  wire n15487_o;
  wire n15488_o;
  wire n15489_o;
  wire n15490_o;
  wire n15492_o;
  wire n15493_o;
  wire [1:0] n15494_o;
  wire n15500_o;
  wire n15501_o;
  wire n15502_o;
  wire n15504_o;
  wire n15506_o;
  wire n15507_o;
  wire n15508_o;
  wire n15509_o;
  wire n15510_o;
  wire n15512_o;
  wire n15513_o;
  wire [1:0] n15514_o;
  wire n15520_o;
  wire n15521_o;
  wire n15522_o;
  wire n15524_o;
  wire n15526_o;
  wire n15527_o;
  wire n15528_o;
  wire n15529_o;
  wire n15530_o;
  wire n15532_o;
  wire n15533_o;
  wire [1:0] n15534_o;
  wire n15540_o;
  wire n15541_o;
  wire n15542_o;
  wire n15544_o;
  wire n15546_o;
  wire n15547_o;
  wire n15548_o;
  wire n15549_o;
  wire n15550_o;
  wire n15552_o;
  wire n15553_o;
  wire [1:0] n15554_o;
  wire n15560_o;
  wire n15561_o;
  wire n15562_o;
  wire n15564_o;
  wire n15566_o;
  wire n15567_o;
  wire n15568_o;
  wire n15569_o;
  wire n15570_o;
  wire n15572_o;
  wire n15577_o;
  wire n15579_o;
  wire n15580_o;
  wire n15581_o;
  wire n15582_o;
  wire n15583_o;
  wire n15584_o;
  wire n15585_o;
  wire n15586_o;
  wire n15589_o;
  wire n15590_o;
  wire n15592_o;
  wire n15593_o;
  wire n15594_o;
  wire n15595_o;
  wire n15596_o;
  wire n15601_o;
  wire n15602_o;
  wire n15603_o;
  wire n15604_o;
  wire n15605_o;
  wire n15607_o;
  wire n15613_o;
  wire n15615_o;
  wire n15618_o;
  wire n15619_o;
  wire n15621_o;
  wire n15622_o;
  wire n15623_o;
  wire n15624_o;
  wire n15625_o;
  wire n15630_o;
  wire n15631_o;
  wire n15632_o;
  wire n15633_o;
  wire n15634_o;
  wire n15636_o;
  wire n15642_o;
  wire n15644_o;
  wire n15647_o;
  wire n15648_o;
  wire n15650_o;
  wire n15651_o;
  wire n15652_o;
  wire n15653_o;
  wire n15654_o;
  wire n15659_o;
  wire n15660_o;
  wire n15661_o;
  wire n15662_o;
  wire n15663_o;
  wire n15665_o;
  wire n15671_o;
  wire n15673_o;
  wire n15676_o;
  wire n15677_o;
  wire n15679_o;
  wire n15680_o;
  wire n15681_o;
  wire n15682_o;
  wire n15683_o;
  wire n15688_o;
  wire n15689_o;
  wire n15690_o;
  wire n15691_o;
  wire n15692_o;
  wire n15694_o;
  wire n15700_o;
  wire n15702_o;
  wire n15705_o;
  wire n15706_o;
  wire n15708_o;
  wire n15709_o;
  wire n15710_o;
  wire n15711_o;
  wire n15712_o;
  wire n15717_o;
  wire n15718_o;
  wire n15719_o;
  wire n15720_o;
  wire n15721_o;
  wire n15723_o;
  wire n15729_o;
  wire n15731_o;
  wire n15734_o;
  wire n15735_o;
  wire n15737_o;
  wire n15738_o;
  wire n15739_o;
  wire n15740_o;
  wire n15741_o;
  wire n15746_o;
  wire n15747_o;
  wire n15748_o;
  wire n15749_o;
  wire n15750_o;
  wire n15752_o;
  wire n15758_o;
  wire n15760_o;
  wire n15763_o;
  wire n15764_o;
  wire n15766_o;
  wire n15767_o;
  wire n15768_o;
  wire n15769_o;
  wire n15770_o;
  wire n15775_o;
  wire n15776_o;
  wire n15777_o;
  wire n15778_o;
  wire n15779_o;
  wire n15781_o;
  wire n15787_o;
  wire n15789_o;
  wire n15792_o;
  wire n15793_o;
  wire n15795_o;
  wire n15796_o;
  wire n15797_o;
  wire n15798_o;
  wire n15799_o;
  wire n15804_o;
  wire n15805_o;
  wire n15806_o;
  wire n15807_o;
  wire n15808_o;
  wire n15810_o;
  wire n15816_o;
  wire n15818_o;
  wire n15821_o;
  wire n15822_o;
  wire n15824_o;
  wire n15825_o;
  wire n15826_o;
  wire n15827_o;
  wire n15828_o;
  wire n15833_o;
  wire n15834_o;
  wire n15835_o;
  wire n15836_o;
  wire n15837_o;
  wire n15839_o;
  wire n15845_o;
  wire n15847_o;
  wire n15850_o;
  wire n15851_o;
  wire n15853_o;
  wire n15854_o;
  wire n15855_o;
  wire n15856_o;
  wire n15857_o;
  wire n15862_o;
  wire n15863_o;
  wire n15864_o;
  wire n15865_o;
  wire n15866_o;
  wire n15868_o;
  wire n15874_o;
  wire n15876_o;
  wire n15879_o;
  wire n15880_o;
  wire n15882_o;
  wire n15883_o;
  wire n15884_o;
  wire n15885_o;
  wire n15886_o;
  wire n15891_o;
  wire n15892_o;
  wire n15893_o;
  wire n15894_o;
  wire n15895_o;
  wire n15897_o;
  wire n15903_o;
  wire n15905_o;
  wire n15908_o;
  wire n15909_o;
  wire n15911_o;
  wire n15912_o;
  wire n15913_o;
  wire n15914_o;
  wire n15915_o;
  wire n15920_o;
  wire n15921_o;
  wire n15922_o;
  wire n15923_o;
  wire n15924_o;
  wire n15926_o;
  wire n15932_o;
  wire n15934_o;
  wire n15936_o;
  wire n15937_o;
  wire n15938_o;
  wire n15939_o;
  wire n15940_o;
  wire n15941_o;
  wire n15942_o;
  wire n15943_o;
  wire n15944_o;
  wire n15945_o;
  wire n15947_o;
  wire n15948_o;
  wire n15953_o;
  wire n15954_o;
  wire n15955_o;
  wire n15957_o;
  wire n15958_o;
  wire n15959_o;
  wire n15964_o;
  wire n15965_o;
  wire n15966_o;
  wire n15967_o;
  wire n15968_o;
  wire n15969_o;
  wire n15970_o;
  wire n15971_o;
  wire n15972_o;
  wire n15975_o;
  wire n15976_o;
  wire n15977_o;
  wire n15978_o;
  wire n15979_o;
  wire n15984_o;
  wire n15985_o;
  wire n15986_o;
  wire n15987_o;
  wire n15988_o;
  wire n15989_o;
  wire n15990_o;
  wire n15993_o;
  wire n15994_o;
  wire n15996_o;
  wire n15997_o;
  wire n15998_o;
  wire n15999_o;
  wire n16000_o;
  wire n16005_o;
  wire n16006_o;
  wire n16007_o;
  wire n16008_o;
  wire n16009_o;
  wire n16010_o;
  wire n16011_o;
  wire n16014_o;
  wire n16015_o;
  wire n16017_o;
  wire n16018_o;
  wire n16019_o;
  wire n16020_o;
  wire n16021_o;
  wire n16026_o;
  wire n16027_o;
  wire n16028_o;
  wire n16029_o;
  wire n16030_o;
  wire n16032_o;
  wire n16033_o;
  wire n16038_o;
  wire n16040_o;
  wire n16041_o;
  wire n16042_o;
  wire n16043_o;
  wire n16044_o;
  wire n16046_o;
  wire n16047_o;
  wire n16048_o;
  wire n16049_o;
  wire n16050_o;
  wire n16055_o;
  wire n16056_o;
  wire n16057_o;
  wire n16058_o;
  wire n16059_o;
  wire n16061_o;
  wire n16062_o;
  wire n16067_o;
  wire n16069_o;
  wire n16071_o;
  wire n16072_o;
  wire n16077_o;
  wire n16079_o;
  wire n16080_o;
  wire n16081_o;
  wire n16083_o;
  wire n16084_o;
  wire n16085_o;
  wire n16086_o;
  wire n16087_o;
  wire n16092_o;
  wire n16093_o;
  wire n16094_o;
  wire n16095_o;
  wire n16096_o;
  wire n16098_o;
  wire n16099_o;
  wire n16104_o;
  wire n16106_o;
  wire n16108_o;
  wire n16109_o;
  wire n16114_o;
  wire n16116_o;
  wire n16117_o;
  wire n16118_o;
  wire n16120_o;
  wire n16121_o;
  wire n16122_o;
  wire n16123_o;
  wire n16124_o;
  wire n16129_o;
  wire n16130_o;
  wire n16131_o;
  wire n16132_o;
  wire n16133_o;
  wire n16135_o;
  wire n16136_o;
  wire n16141_o;
  wire n16143_o;
  wire n16145_o;
  wire n16146_o;
  wire n16151_o;
  wire n16153_o;
  wire n16154_o;
  wire n16155_o;
  wire n16157_o;
  wire n16158_o;
  wire n16159_o;
  wire n16160_o;
  wire n16161_o;
  wire n16166_o;
  wire n16167_o;
  wire n16168_o;
  wire n16169_o;
  wire n16170_o;
  wire n16172_o;
  wire n16173_o;
  wire n16178_o;
  wire n16180_o;
  wire n16182_o;
  wire n16183_o;
  wire n16188_o;
  wire n16190_o;
  wire n16191_o;
  wire n16192_o;
  wire n16194_o;
  wire n16195_o;
  wire n16196_o;
  wire n16197_o;
  wire n16198_o;
  wire n16203_o;
  wire n16204_o;
  wire n16205_o;
  wire n16206_o;
  wire n16207_o;
  wire n16209_o;
  wire n16210_o;
  wire n16215_o;
  wire n16217_o;
  wire n16219_o;
  wire n16220_o;
  wire n16225_o;
  wire n16227_o;
  wire n16228_o;
  wire n16229_o;
  wire n16231_o;
  wire n16232_o;
  wire n16233_o;
  wire n16234_o;
  wire n16235_o;
  wire n16240_o;
  wire n16241_o;
  wire n16242_o;
  wire n16243_o;
  wire n16244_o;
  wire n16246_o;
  wire n16247_o;
  wire n16252_o;
  wire n16254_o;
  wire n16256_o;
  wire n16257_o;
  wire n16262_o;
  wire n16264_o;
  wire n16265_o;
  wire n16266_o;
  wire n16268_o;
  wire n16269_o;
  wire n16270_o;
  wire n16271_o;
  wire n16272_o;
  wire n16277_o;
  wire n16278_o;
  wire n16279_o;
  wire n16280_o;
  wire n16281_o;
  wire n16283_o;
  wire n16284_o;
  wire n16289_o;
  wire n16291_o;
  wire n16293_o;
  wire n16294_o;
  wire n16299_o;
  wire n16301_o;
  wire n16302_o;
  wire n16303_o;
  wire n16305_o;
  wire n16306_o;
  wire n16307_o;
  wire n16308_o;
  wire n16309_o;
  wire n16314_o;
  wire n16315_o;
  wire n16316_o;
  wire n16317_o;
  wire n16318_o;
  wire n16320_o;
  wire n16321_o;
  wire n16326_o;
  wire n16328_o;
  wire n16330_o;
  wire n16331_o;
  wire n16336_o;
  wire n16338_o;
  wire n16339_o;
  wire n16340_o;
  wire n16342_o;
  wire n16343_o;
  wire n16344_o;
  wire n16345_o;
  wire n16346_o;
  wire n16351_o;
  wire n16352_o;
  wire n16353_o;
  wire n16354_o;
  wire n16355_o;
  wire n16357_o;
  wire n16358_o;
  wire n16363_o;
  wire n16365_o;
  wire n16367_o;
  wire n16368_o;
  wire n16373_o;
  wire n16375_o;
  wire n16376_o;
  wire n16377_o;
  wire n16379_o;
  wire n16380_o;
  wire n16381_o;
  wire n16382_o;
  wire n16383_o;
  wire n16388_o;
  wire n16389_o;
  wire n16390_o;
  wire n16391_o;
  wire n16392_o;
  wire n16394_o;
  wire n16395_o;
  wire n16400_o;
  wire n16402_o;
  wire n16404_o;
  wire n16405_o;
  wire n16410_o;
  wire n16412_o;
  wire n16413_o;
  wire n16414_o;
  wire n16416_o;
  wire n16417_o;
  wire n16418_o;
  wire n16419_o;
  wire n16424_o;
  wire n16425_o;
  wire n16426_o;
  wire n16427_o;
  wire n16429_o;
  wire n16430_o;
  wire n16431_o;
  wire n16436_o;
  wire n16437_o;
  wire n16438_o;
  wire n16439_o;
  wire n16441_o;
  wire n16442_o;
  wire n16447_o;
  wire n16448_o;
  wire n16449_o;
  wire n16451_o;
  wire n16452_o;
  wire n16453_o;
  wire n16458_o;
  wire n16459_o;
  wire n16460_o;
  wire n16461_o;
  wire n16462_o;
  wire n16463_o;
  wire n16464_o;
  wire n16465_o;
  wire n16466_o;
  wire n16469_o;
  wire n16470_o;
  wire n16471_o;
  wire n16472_o;
  wire n16473_o;
  wire n16478_o;
  wire n16479_o;
  wire n16480_o;
  wire n16481_o;
  wire n16482_o;
  wire n16483_o;
  wire n16484_o;
  wire n16487_o;
  wire n16488_o;
  wire n16490_o;
  wire n16491_o;
  wire n16492_o;
  wire n16493_o;
  wire n16494_o;
  wire n16499_o;
  wire n16500_o;
  wire n16501_o;
  wire n16502_o;
  wire n16503_o;
  wire n16504_o;
  wire n16505_o;
  wire n16508_o;
  wire n16509_o;
  wire n16511_o;
  wire n16512_o;
  wire n16513_o;
  wire n16514_o;
  wire n16515_o;
  wire n16520_o;
  wire n16521_o;
  wire n16522_o;
  wire n16523_o;
  wire n16524_o;
  wire n16526_o;
  wire n16527_o;
  wire n16528_o;
  wire n16533_o;
  wire n16534_o;
  wire n16536_o;
  wire n16537_o;
  wire n16538_o;
  wire n16543_o;
  wire n16544_o;
  wire n16545_o;
  wire n16546_o;
  wire n16548_o;
  wire n16549_o;
  wire n16550_o;
  wire n16551_o;
  wire n16552_o;
  wire n16557_o;
  wire n16558_o;
  wire n16559_o;
  wire n16560_o;
  wire n16561_o;
  wire n16563_o;
  wire n16564_o;
  wire n16565_o;
  wire n16570_o;
  wire n16571_o;
  wire n16573_o;
  wire n16574_o;
  wire n16575_o;
  wire n16580_o;
  wire n16581_o;
  wire n16582_o;
  wire n16583_o;
  wire n16585_o;
  wire n16586_o;
  wire n16587_o;
  wire n16588_o;
  wire n16589_o;
  wire n16594_o;
  wire n16595_o;
  wire n16596_o;
  wire n16597_o;
  wire n16598_o;
  wire n16600_o;
  wire n16601_o;
  wire n16602_o;
  wire n16607_o;
  wire n16608_o;
  wire n16610_o;
  wire n16611_o;
  wire n16612_o;
  wire n16617_o;
  wire n16618_o;
  wire n16619_o;
  wire n16620_o;
  wire n16622_o;
  wire n16623_o;
  wire n16624_o;
  wire n16625_o;
  wire n16626_o;
  wire n16631_o;
  wire n16632_o;
  wire n16633_o;
  wire n16634_o;
  wire n16635_o;
  wire n16637_o;
  wire n16638_o;
  wire n16639_o;
  wire n16644_o;
  wire n16645_o;
  wire n16647_o;
  wire n16648_o;
  wire n16649_o;
  wire n16654_o;
  wire n16655_o;
  wire n16656_o;
  wire n16657_o;
  wire n16659_o;
  wire n16660_o;
  wire n16661_o;
  wire n16662_o;
  wire n16663_o;
  wire n16668_o;
  wire n16669_o;
  wire n16670_o;
  wire n16671_o;
  wire n16672_o;
  wire n16674_o;
  wire n16675_o;
  wire n16676_o;
  wire n16681_o;
  wire n16682_o;
  wire n16684_o;
  wire n16685_o;
  wire n16686_o;
  wire n16691_o;
  wire n16692_o;
  wire n16693_o;
  wire n16694_o;
  wire n16696_o;
  wire n16697_o;
  wire n16698_o;
  wire n16699_o;
  wire n16700_o;
  wire n16705_o;
  wire n16706_o;
  wire n16707_o;
  wire n16708_o;
  wire n16709_o;
  wire n16711_o;
  wire n16712_o;
  wire n16713_o;
  wire n16718_o;
  wire n16719_o;
  wire n16721_o;
  wire n16722_o;
  wire n16723_o;
  wire n16728_o;
  wire n16729_o;
  wire n16730_o;
  wire n16731_o;
  wire n16733_o;
  wire n16734_o;
  wire n16735_o;
  wire n16736_o;
  wire n16737_o;
  wire n16742_o;
  wire n16743_o;
  wire n16744_o;
  wire n16745_o;
  wire n16746_o;
  wire n16748_o;
  wire n16749_o;
  wire n16750_o;
  wire n16755_o;
  wire n16756_o;
  wire n16758_o;
  wire n16759_o;
  wire n16760_o;
  wire n16765_o;
  wire n16766_o;
  wire n16767_o;
  wire n16768_o;
  wire n16770_o;
  wire n16771_o;
  wire n16772_o;
  wire n16773_o;
  wire n16774_o;
  wire n16779_o;
  wire n16780_o;
  wire n16781_o;
  wire n16782_o;
  wire n16783_o;
  wire n16785_o;
  wire n16786_o;
  wire n16787_o;
  wire n16792_o;
  wire n16793_o;
  wire n16795_o;
  wire n16796_o;
  wire n16797_o;
  wire n16802_o;
  wire n16803_o;
  wire n16804_o;
  wire n16805_o;
  wire n16807_o;
  wire n16808_o;
  wire n16809_o;
  wire n16810_o;
  wire n16811_o;
  wire n16816_o;
  wire n16817_o;
  wire n16818_o;
  wire n16819_o;
  wire n16820_o;
  wire n16822_o;
  wire n16823_o;
  wire n16824_o;
  wire n16829_o;
  wire n16830_o;
  wire n16832_o;
  wire n16833_o;
  wire n16834_o;
  wire n16839_o;
  wire n16840_o;
  wire n16841_o;
  wire n16842_o;
  wire n16844_o;
  wire n16845_o;
  wire n16846_o;
  wire n16847_o;
  wire n16848_o;
  wire n16853_o;
  wire n16854_o;
  wire n16855_o;
  wire n16856_o;
  wire n16857_o;
  wire n16859_o;
  wire n16860_o;
  wire n16861_o;
  wire n16866_o;
  wire n16867_o;
  wire n16869_o;
  wire n16870_o;
  wire n16871_o;
  wire n16876_o;
  wire n16877_o;
  wire n16878_o;
  wire n16879_o;
  wire n16881_o;
  wire n16882_o;
  wire n16883_o;
  wire n16884_o;
  wire n16885_o;
  wire n16890_o;
  wire n16891_o;
  wire n16892_o;
  wire n16893_o;
  wire n16894_o;
  wire n16896_o;
  wire n16897_o;
  wire n16898_o;
  wire n16903_o;
  wire n16904_o;
  wire n16906_o;
  wire n16907_o;
  wire n16908_o;
  wire n16913_o;
  wire n16914_o;
  wire n16915_o;
  wire n16916_o;
  wire n16918_o;
  wire n16919_o;
  wire n16920_o;
  wire n16921_o;
  wire n16926_o;
  wire n16927_o;
  wire n16928_o;
  wire n16929_o;
  wire n16931_o;
  wire n16932_o;
  wire n16933_o;
  wire n16938_o;
  wire n16939_o;
  wire n16940_o;
  wire n16941_o;
  wire n16943_o;
  wire n16944_o;
  wire n16949_o;
  wire n16950_o;
  wire n16951_o;
  wire n16953_o;
  wire n16954_o;
  wire n16955_o;
  wire n16960_o;
  wire n16961_o;
  wire n16962_o;
  wire n16963_o;
  wire n16964_o;
  wire n16965_o;
  wire n16966_o;
  wire n16967_o;
  wire n16968_o;
  wire n16971_o;
  wire n16972_o;
  wire n16973_o;
  wire n16974_o;
  wire n16975_o;
  wire n16980_o;
  wire n16981_o;
  wire n16982_o;
  wire n16983_o;
  wire n16984_o;
  wire n16985_o;
  wire n16986_o;
  wire n16989_o;
  wire n16990_o;
  wire n16992_o;
  wire n16993_o;
  wire n16994_o;
  wire n16995_o;
  wire n16996_o;
  wire n17001_o;
  wire n17002_o;
  wire n17003_o;
  wire n17004_o;
  wire n17005_o;
  wire n17006_o;
  wire n17007_o;
  wire n17010_o;
  wire n17011_o;
  wire n17013_o;
  wire n17014_o;
  wire n17015_o;
  wire n17016_o;
  wire n17017_o;
  wire n17022_o;
  wire n17023_o;
  wire n17024_o;
  wire n17025_o;
  wire n17026_o;
  wire n17028_o;
  wire n17029_o;
  wire n17030_o;
  wire n17035_o;
  wire n17036_o;
  wire n17038_o;
  wire n17039_o;
  wire n17040_o;
  wire n17045_o;
  wire n17046_o;
  wire n17047_o;
  wire n17048_o;
  wire n17050_o;
  wire n17051_o;
  wire n17052_o;
  wire n17053_o;
  wire n17054_o;
  wire n17059_o;
  wire n17060_o;
  wire n17061_o;
  wire n17062_o;
  wire n17063_o;
  wire n17065_o;
  wire n17066_o;
  wire n17067_o;
  wire n17072_o;
  wire n17073_o;
  wire n17075_o;
  wire n17076_o;
  wire n17077_o;
  wire n17082_o;
  wire n17083_o;
  wire n17084_o;
  wire n17085_o;
  wire n17087_o;
  wire n17088_o;
  wire n17089_o;
  wire n17090_o;
  wire n17091_o;
  wire n17096_o;
  wire n17097_o;
  wire n17098_o;
  wire n17099_o;
  wire n17100_o;
  wire n17102_o;
  wire n17103_o;
  wire n17104_o;
  wire n17109_o;
  wire n17110_o;
  wire n17112_o;
  wire n17113_o;
  wire n17114_o;
  wire n17119_o;
  wire n17120_o;
  wire n17121_o;
  wire n17122_o;
  wire n17124_o;
  wire n17125_o;
  wire n17126_o;
  wire n17127_o;
  wire n17128_o;
  wire n17133_o;
  wire n17134_o;
  wire n17135_o;
  wire n17136_o;
  wire n17137_o;
  wire n17139_o;
  wire n17140_o;
  wire n17141_o;
  wire n17146_o;
  wire n17147_o;
  wire n17149_o;
  wire n17150_o;
  wire n17151_o;
  wire n17156_o;
  wire n17157_o;
  wire n17158_o;
  wire n17159_o;
  wire n17161_o;
  wire n17162_o;
  wire n17163_o;
  wire n17164_o;
  wire n17165_o;
  wire n17170_o;
  wire n17171_o;
  wire n17172_o;
  wire n17173_o;
  wire n17174_o;
  wire n17176_o;
  wire n17177_o;
  wire n17178_o;
  wire n17183_o;
  wire n17184_o;
  wire n17186_o;
  wire n17187_o;
  wire n17188_o;
  wire n17193_o;
  wire n17194_o;
  wire n17195_o;
  wire n17196_o;
  wire n17198_o;
  wire n17199_o;
  wire n17200_o;
  wire n17201_o;
  wire n17202_o;
  wire n17207_o;
  wire n17208_o;
  wire n17209_o;
  wire n17210_o;
  wire n17211_o;
  wire n17213_o;
  wire n17214_o;
  wire n17215_o;
  wire n17220_o;
  wire n17221_o;
  wire n17223_o;
  wire n17224_o;
  wire n17225_o;
  wire n17230_o;
  wire n17231_o;
  wire n17232_o;
  wire n17233_o;
  wire n17235_o;
  wire n17236_o;
  wire n17237_o;
  wire n17238_o;
  wire n17239_o;
  wire n17244_o;
  wire n17245_o;
  wire n17246_o;
  wire n17247_o;
  wire n17248_o;
  wire n17250_o;
  wire n17251_o;
  wire n17252_o;
  wire n17257_o;
  wire n17258_o;
  wire n17260_o;
  wire n17261_o;
  wire n17262_o;
  wire n17267_o;
  wire n17268_o;
  wire n17269_o;
  wire n17270_o;
  wire n17272_o;
  wire n17273_o;
  wire n17274_o;
  wire n17275_o;
  wire n17276_o;
  wire n17281_o;
  wire n17282_o;
  wire n17283_o;
  wire n17284_o;
  wire n17285_o;
  wire n17287_o;
  wire n17288_o;
  wire n17289_o;
  wire n17294_o;
  wire n17295_o;
  wire n17297_o;
  wire n17298_o;
  wire n17299_o;
  wire n17304_o;
  wire n17305_o;
  wire n17306_o;
  wire n17307_o;
  wire n17309_o;
  wire n17310_o;
  wire n17311_o;
  wire n17312_o;
  wire n17313_o;
  wire n17318_o;
  wire n17319_o;
  wire n17320_o;
  wire n17321_o;
  wire n17322_o;
  wire n17324_o;
  wire n17325_o;
  wire n17326_o;
  wire n17331_o;
  wire n17332_o;
  wire n17334_o;
  wire n17335_o;
  wire n17336_o;
  wire n17341_o;
  wire n17342_o;
  wire n17343_o;
  wire n17344_o;
  wire n17346_o;
  wire n17347_o;
  wire n17348_o;
  wire n17349_o;
  wire n17350_o;
  wire n17355_o;
  wire n17356_o;
  wire n17357_o;
  wire n17358_o;
  wire n17359_o;
  wire n17361_o;
  wire n17362_o;
  wire n17363_o;
  wire n17368_o;
  wire n17369_o;
  wire n17371_o;
  wire n17372_o;
  wire n17373_o;
  wire n17378_o;
  wire n17379_o;
  wire n17380_o;
  wire n17381_o;
  wire n17383_o;
  wire n17384_o;
  wire n17385_o;
  wire n17386_o;
  wire n17387_o;
  wire n17392_o;
  wire n17393_o;
  wire n17394_o;
  wire n17395_o;
  wire n17396_o;
  wire n17398_o;
  wire n17399_o;
  wire n17400_o;
  wire n17405_o;
  wire n17406_o;
  wire n17408_o;
  wire n17409_o;
  wire n17410_o;
  wire n17415_o;
  wire n17416_o;
  wire n17417_o;
  wire n17418_o;
  wire n17420_o;
  wire n17421_o;
  wire n17422_o;
  wire n17423_o;
  wire n17428_o;
  wire n17429_o;
  wire n17430_o;
  wire n17431_o;
  wire n17433_o;
  wire n17434_o;
  wire n17435_o;
  wire n17440_o;
  wire n17441_o;
  wire n17442_o;
  wire n17443_o;
  wire n17445_o;
  wire n17446_o;
  wire n17451_o;
  wire n17452_o;
  wire n17453_o;
  wire n17455_o;
  wire n17456_o;
  wire n17457_o;
  wire n17462_o;
  wire n17463_o;
  wire n17464_o;
  wire n17465_o;
  wire n17466_o;
  wire n17467_o;
  wire n17468_o;
  wire n17469_o;
  wire n17470_o;
  wire n17473_o;
  wire n17474_o;
  wire n17475_o;
  wire n17476_o;
  wire n17477_o;
  wire n17482_o;
  wire n17483_o;
  wire n17484_o;
  wire n17485_o;
  wire n17486_o;
  wire n17487_o;
  wire n17488_o;
  wire n17491_o;
  wire n17492_o;
  wire n17494_o;
  wire n17495_o;
  wire n17496_o;
  wire n17497_o;
  wire n17498_o;
  wire n17503_o;
  wire n17504_o;
  wire n17505_o;
  wire n17506_o;
  wire n17507_o;
  wire n17508_o;
  wire n17509_o;
  wire n17512_o;
  wire n17513_o;
  wire n17515_o;
  wire n17516_o;
  wire n17517_o;
  wire n17518_o;
  wire n17519_o;
  wire n17524_o;
  wire n17525_o;
  wire n17526_o;
  wire n17527_o;
  wire n17528_o;
  wire n17530_o;
  wire n17531_o;
  wire n17532_o;
  wire n17537_o;
  wire n17538_o;
  wire n17540_o;
  wire n17541_o;
  wire n17542_o;
  wire n17547_o;
  wire n17548_o;
  wire n17549_o;
  wire n17550_o;
  wire n17552_o;
  wire n17553_o;
  wire n17554_o;
  wire n17555_o;
  wire n17556_o;
  wire n17561_o;
  wire n17562_o;
  wire n17563_o;
  wire n17564_o;
  wire n17565_o;
  wire n17567_o;
  wire n17568_o;
  wire n17569_o;
  wire n17574_o;
  wire n17575_o;
  wire n17577_o;
  wire n17578_o;
  wire n17579_o;
  wire n17584_o;
  wire n17585_o;
  wire n17586_o;
  wire n17587_o;
  wire n17589_o;
  wire n17590_o;
  wire n17591_o;
  wire n17592_o;
  wire n17593_o;
  wire n17598_o;
  wire n17599_o;
  wire n17600_o;
  wire n17601_o;
  wire n17602_o;
  wire n17604_o;
  wire n17605_o;
  wire n17606_o;
  wire n17611_o;
  wire n17612_o;
  wire n17614_o;
  wire n17615_o;
  wire n17616_o;
  wire n17621_o;
  wire n17622_o;
  wire n17623_o;
  wire n17624_o;
  wire n17626_o;
  wire n17627_o;
  wire n17628_o;
  wire n17629_o;
  wire n17630_o;
  wire n17635_o;
  wire n17636_o;
  wire n17637_o;
  wire n17638_o;
  wire n17639_o;
  wire n17641_o;
  wire n17642_o;
  wire n17643_o;
  wire n17648_o;
  wire n17649_o;
  wire n17651_o;
  wire n17652_o;
  wire n17653_o;
  wire n17658_o;
  wire n17659_o;
  wire n17660_o;
  wire n17661_o;
  wire n17663_o;
  wire n17664_o;
  wire n17665_o;
  wire n17666_o;
  wire n17667_o;
  wire n17672_o;
  wire n17673_o;
  wire n17674_o;
  wire n17675_o;
  wire n17676_o;
  wire n17678_o;
  wire n17679_o;
  wire n17680_o;
  wire n17685_o;
  wire n17686_o;
  wire n17688_o;
  wire n17689_o;
  wire n17690_o;
  wire n17695_o;
  wire n17696_o;
  wire n17697_o;
  wire n17698_o;
  wire n17700_o;
  wire n17701_o;
  wire n17702_o;
  wire n17703_o;
  wire n17704_o;
  wire n17709_o;
  wire n17710_o;
  wire n17711_o;
  wire n17712_o;
  wire n17713_o;
  wire n17715_o;
  wire n17716_o;
  wire n17717_o;
  wire n17722_o;
  wire n17723_o;
  wire n17725_o;
  wire n17726_o;
  wire n17727_o;
  wire n17732_o;
  wire n17733_o;
  wire n17734_o;
  wire n17735_o;
  wire n17737_o;
  wire n17738_o;
  wire n17739_o;
  wire n17740_o;
  wire n17741_o;
  wire n17746_o;
  wire n17747_o;
  wire n17748_o;
  wire n17749_o;
  wire n17750_o;
  wire n17752_o;
  wire n17753_o;
  wire n17754_o;
  wire n17759_o;
  wire n17760_o;
  wire n17762_o;
  wire n17763_o;
  wire n17764_o;
  wire n17769_o;
  wire n17770_o;
  wire n17771_o;
  wire n17772_o;
  wire n17774_o;
  wire n17775_o;
  wire n17776_o;
  wire n17777_o;
  wire n17778_o;
  wire n17783_o;
  wire n17784_o;
  wire n17785_o;
  wire n17786_o;
  wire n17787_o;
  wire n17789_o;
  wire n17790_o;
  wire n17791_o;
  wire n17796_o;
  wire n17797_o;
  wire n17799_o;
  wire n17800_o;
  wire n17801_o;
  wire n17806_o;
  wire n17807_o;
  wire n17808_o;
  wire n17809_o;
  wire n17811_o;
  wire n17812_o;
  wire n17813_o;
  wire n17814_o;
  wire n17815_o;
  wire n17820_o;
  wire n17821_o;
  wire n17822_o;
  wire n17823_o;
  wire n17824_o;
  wire n17826_o;
  wire n17827_o;
  wire n17828_o;
  wire n17833_o;
  wire n17834_o;
  wire n17836_o;
  wire n17837_o;
  wire n17838_o;
  wire n17843_o;
  wire n17844_o;
  wire n17845_o;
  wire n17846_o;
  wire n17848_o;
  wire n17849_o;
  wire n17850_o;
  wire n17851_o;
  wire n17852_o;
  wire n17857_o;
  wire n17858_o;
  wire n17859_o;
  wire n17860_o;
  wire n17861_o;
  wire n17863_o;
  wire n17864_o;
  wire n17865_o;
  wire n17870_o;
  wire n17871_o;
  wire n17873_o;
  wire n17874_o;
  wire n17875_o;
  wire n17880_o;
  wire n17881_o;
  wire n17882_o;
  wire n17883_o;
  wire n17885_o;
  wire n17886_o;
  wire n17887_o;
  wire n17888_o;
  wire n17889_o;
  wire n17894_o;
  wire n17895_o;
  wire n17896_o;
  wire n17897_o;
  wire n17898_o;
  wire n17900_o;
  wire n17901_o;
  wire n17902_o;
  wire n17907_o;
  wire n17908_o;
  wire n17910_o;
  wire n17911_o;
  wire n17912_o;
  wire n17917_o;
  wire n17918_o;
  wire n17919_o;
  wire n17920_o;
  wire n17922_o;
  wire n17923_o;
  wire n17924_o;
  wire n17925_o;
  wire n17930_o;
  wire n17931_o;
  wire n17932_o;
  wire n17933_o;
  wire n17934_o;
  wire n17941_o;
  wire n17943_o;
  wire [11:0] n17945_o;
  wire n17948_o;
  wire n17954_o;
  wire n17955_o;
  wire n17956_o;
  wire n17957_o;
  wire n17958_o;
  wire n17959_o;
  wire n17960_o;
  wire n17961_o;
  wire n17962_o;
  wire n17963_o;
  wire n17964_o;
  wire n17970_o;
  wire n17971_o;
  wire n17972_o;
  wire n17973_o;
  wire n17974_o;
  wire n17975_o;
  wire n17976_o;
  wire n17977_o;
  wire n17978_o;
  wire n17979_o;
  wire n17980_o;
  wire n17986_o;
  wire n17987_o;
  wire n17988_o;
  wire n17989_o;
  wire n17990_o;
  wire n17991_o;
  wire n17992_o;
  wire n17993_o;
  wire n17994_o;
  wire n17995_o;
  wire n17996_o;
  wire n18002_o;
  wire n18003_o;
  wire n18004_o;
  wire n18005_o;
  wire n18006_o;
  wire n18007_o;
  wire n18008_o;
  wire n18009_o;
  wire n18010_o;
  wire n18011_o;
  wire n18012_o;
  wire n18018_o;
  wire n18019_o;
  wire n18020_o;
  wire n18021_o;
  wire n18022_o;
  wire n18023_o;
  wire n18024_o;
  wire n18025_o;
  wire n18026_o;
  wire n18027_o;
  wire n18028_o;
  wire n18034_o;
  wire n18035_o;
  wire n18036_o;
  wire n18037_o;
  wire n18038_o;
  wire n18039_o;
  wire n18040_o;
  wire n18041_o;
  wire n18042_o;
  wire n18043_o;
  wire n18044_o;
  wire n18050_o;
  wire n18051_o;
  wire n18052_o;
  wire n18053_o;
  wire n18054_o;
  wire n18055_o;
  wire n18056_o;
  wire n18057_o;
  wire n18058_o;
  wire n18059_o;
  wire n18060_o;
  wire n18066_o;
  wire n18067_o;
  wire n18068_o;
  wire n18069_o;
  wire n18070_o;
  wire n18071_o;
  wire n18072_o;
  wire n18073_o;
  wire n18074_o;
  wire n18075_o;
  wire n18076_o;
  wire n18082_o;
  wire n18083_o;
  wire n18084_o;
  wire n18085_o;
  wire n18086_o;
  wire n18087_o;
  wire n18088_o;
  wire n18089_o;
  wire n18090_o;
  wire n18091_o;
  wire n18092_o;
  wire n18098_o;
  wire n18099_o;
  wire n18100_o;
  wire n18101_o;
  wire n18102_o;
  wire n18103_o;
  wire n18104_o;
  wire n18105_o;
  wire n18106_o;
  wire n18107_o;
  wire n18108_o;
  wire n18114_o;
  wire n18115_o;
  wire n18116_o;
  wire n18117_o;
  wire n18118_o;
  wire n18119_o;
  wire n18120_o;
  wire n18121_o;
  wire n18122_o;
  wire n18123_o;
  wire n18124_o;
  wire n18130_o;
  wire n18131_o;
  wire n18132_o;
  wire n18133_o;
  wire n18134_o;
  wire n18135_o;
  wire n18136_o;
  wire n18137_o;
  wire n18138_o;
  wire n18139_o;
  wire n18140_o;
  wire n18141_o;
  wire n18147_o;
  wire n18148_o;
  wire n18149_o;
  wire n18156_o;
  wire n18158_o;
  wire n18162_o;
  wire n18166_o;
  wire n18167_o;
  wire n18173_o;
  wire n18174_o;
  wire n18175_o;
  wire n18177_o;
  wire n18178_o;
  wire n18179_o;
  wire n18184_o;
  wire n18185_o;
  wire n18186_o;
  wire n18187_o;
  wire n18189_o;
  wire n18190_o;
  wire n18191_o;
  wire n18196_o;
  wire n18197_o;
  wire n18204_o;
  wire n18206_o;
  wire n18210_o;
  wire n18214_o;
  wire n18215_o;
  wire n18221_o;
  wire n18222_o;
  wire n18223_o;
  wire n18225_o;
  wire n18226_o;
  wire n18227_o;
  wire n18232_o;
  wire n18233_o;
  wire n18234_o;
  wire n18235_o;
  wire n18237_o;
  wire n18238_o;
  wire n18239_o;
  wire n18244_o;
  wire n18245_o;
  wire n18252_o;
  wire n18254_o;
  wire n18258_o;
  wire n18262_o;
  wire n18263_o;
  wire n18269_o;
  wire n18270_o;
  wire n18271_o;
  wire n18273_o;
  wire n18274_o;
  wire n18275_o;
  wire n18280_o;
  wire n18281_o;
  wire n18282_o;
  wire n18283_o;
  wire n18285_o;
  wire n18286_o;
  wire n18287_o;
  wire n18292_o;
  wire n18293_o;
  wire n18300_o;
  wire n18302_o;
  wire n18306_o;
  wire n18310_o;
  wire n18311_o;
  wire n18317_o;
  wire n18318_o;
  wire n18319_o;
  wire n18321_o;
  wire n18322_o;
  wire n18323_o;
  wire n18328_o;
  wire n18329_o;
  wire n18330_o;
  wire n18331_o;
  wire n18333_o;
  wire n18334_o;
  wire n18335_o;
  wire n18340_o;
  wire n18341_o;
  wire n18348_o;
  wire n18350_o;
  wire n18354_o;
  wire n18358_o;
  wire n18359_o;
  wire n18365_o;
  wire n18366_o;
  wire n18367_o;
  wire n18369_o;
  wire n18370_o;
  wire n18371_o;
  wire n18376_o;
  wire n18377_o;
  wire n18378_o;
  wire n18379_o;
  wire n18381_o;
  wire n18382_o;
  wire n18383_o;
  wire n18388_o;
  wire n18389_o;
  wire n18396_o;
  wire n18398_o;
  wire n18402_o;
  wire n18406_o;
  wire n18407_o;
  wire n18413_o;
  wire n18414_o;
  wire n18415_o;
  wire n18417_o;
  wire n18418_o;
  wire n18419_o;
  wire n18424_o;
  wire n18425_o;
  wire n18426_o;
  wire n18427_o;
  wire n18429_o;
  wire n18430_o;
  wire n18431_o;
  wire n18436_o;
  wire n18437_o;
  wire n18444_o;
  wire n18446_o;
  wire n18450_o;
  wire n18454_o;
  wire n18455_o;
  wire n18461_o;
  wire n18462_o;
  wire n18463_o;
  wire n18465_o;
  wire n18466_o;
  wire n18467_o;
  wire n18472_o;
  wire n18473_o;
  wire n18474_o;
  wire n18475_o;
  wire n18477_o;
  wire n18478_o;
  wire n18479_o;
  wire n18484_o;
  wire n18485_o;
  wire n18492_o;
  wire n18494_o;
  wire n18498_o;
  wire n18502_o;
  wire n18503_o;
  wire n18509_o;
  wire n18510_o;
  wire n18511_o;
  wire n18513_o;
  wire n18514_o;
  wire n18515_o;
  wire n18520_o;
  wire n18521_o;
  wire n18522_o;
  wire n18523_o;
  wire n18525_o;
  wire n18526_o;
  wire n18527_o;
  wire n18532_o;
  wire n18533_o;
  wire n18540_o;
  wire n18542_o;
  wire n18546_o;
  wire n18550_o;
  wire n18551_o;
  wire n18557_o;
  wire n18558_o;
  wire n18559_o;
  wire n18561_o;
  wire n18562_o;
  wire n18563_o;
  wire n18568_o;
  wire n18569_o;
  wire n18570_o;
  wire n18571_o;
  wire n18573_o;
  wire n18574_o;
  wire n18575_o;
  wire n18580_o;
  wire n18581_o;
  wire n18588_o;
  wire n18590_o;
  wire n18594_o;
  wire n18598_o;
  wire n18599_o;
  wire n18605_o;
  wire n18606_o;
  wire n18607_o;
  wire n18609_o;
  wire n18610_o;
  wire n18611_o;
  wire n18616_o;
  wire n18617_o;
  wire n18618_o;
  wire n18619_o;
  wire n18621_o;
  wire n18622_o;
  wire n18623_o;
  wire n18628_o;
  wire n18629_o;
  wire n18636_o;
  wire n18638_o;
  wire n18642_o;
  wire n18646_o;
  wire n18647_o;
  wire n18653_o;
  wire n18654_o;
  wire n18655_o;
  wire n18657_o;
  wire n18658_o;
  wire n18659_o;
  wire n18664_o;
  wire n18665_o;
  wire n18666_o;
  wire n18667_o;
  wire n18669_o;
  wire n18670_o;
  wire n18671_o;
  wire n18676_o;
  wire n18677_o;
  wire n18684_o;
  wire n18686_o;
  wire n18690_o;
  wire n18694_o;
  wire n18695_o;
  wire n18701_o;
  wire n18702_o;
  wire n18703_o;
  wire n18705_o;
  wire n18706_o;
  wire n18707_o;
  wire n18712_o;
  wire n18713_o;
  wire n18714_o;
  wire n18715_o;
  wire n18717_o;
  wire n18718_o;
  wire n18719_o;
  wire n18724_o;
  wire n18725_o;
  wire [11:0] n18726_o;
  wire n18728_o;
  wire n18729_o;
  wire n18730_o;
  wire n18731_o;
  wire n18732_o;
  wire n18737_o;
  wire n18738_o;
  wire [11:0] n18739_o;
  wire n18742_o;
  wire n18743_o;
  wire n18744_o;
  wire n18745_o;
  wire n18750_o;
  wire n18751_o;
  wire n18752_o;
  wire [11:0] n18753_o;
  wire n18756_o;
  wire n18757_o;
  wire n18758_o;
  wire n18759_o;
  wire n18764_o;
  wire n18765_o;
  wire n18766_o;
  wire [11:0] n18767_o;
  wire n18771_o;
  wire n18774_o;
  wire n18777_o;
  wire n18780_o;
  wire n18783_o;
  wire n18786_o;
  wire n18789_o;
  wire n18792_o;
  wire n18795_o;
  wire n18798_o;
  wire n18801_o;
  wire n18804_o;
  wire n18807_o;
  wire n18812_o;
  wire n18813_o;
  wire n18814_o;
  wire n18815_o;
  wire n18816_o;
  wire n18817_o;
  wire n18818_o;
  wire [3:0] n18819_o;
  wire n18821_o;
  wire n18822_o;
  wire n18827_o;
  wire n18828_o;
  wire n18829_o;
  wire n18830_o;
  wire n18831_o;
  wire n18832_o;
  wire n18833_o;
  wire [3:0] n18834_o;
  wire n18839_o;
  wire n18840_o;
  wire n18841_o;
  wire n18842_o;
  wire n18843_o;
  wire n18844_o;
  wire n18845_o;
  wire n18846_o;
  wire n18847_o;
  wire n18848_o;
  wire n18849_o;
  wire n18850_o;
  wire n18851_o;
  wire n18852_o;
  wire n18853_o;
  wire n18854_o;
  wire n18855_o;
  wire n18856_o;
  wire n18857_o;
  wire n18858_o;
  wire n18859_o;
  wire n18860_o;
  wire n18861_o;
  wire n18862_o;
  wire n18863_o;
  wire n18864_o;
  wire n18865_o;
  wire n18866_o;
  wire [3:0] n18867_o;
  wire n18869_o;
  wire n18870_o;
  wire n18875_o;
  wire n18876_o;
  wire n18877_o;
  wire n18879_o;
  wire n18884_o;
  wire n18885_o;
  wire n18886_o;
  wire n18887_o;
  wire n18888_o;
  wire n18889_o;
  wire n18890_o;
  wire [3:0] n18891_o;
  wire n18892_o;
  wire n18899_o;
  wire n18901_o;
  wire [11:0] n18903_o;
  wire [11:0] n18906_o;
  wire [57:0] n18910_o;
  wire [57:0] n18911_o;
  wire [57:0] n18912_o;
  wire [57:0] n18913_o;
  wire [57:0] n18914_o;
  wire [11:0] n18917_o;
  reg [11:0] n18918_q;
  wire [23:0] n18919_o;
  wire n18920_o;
  wire n18921_o;
  reg n18922_q;
  wire n18923_o;
  wire n18924_o;
  reg n18925_q;
  wire n18926_o;
  wire n18927_o;
  reg n18928_q;
  wire n18929_o;
  wire n18930_o;
  reg n18931_q;
  wire n18932_o;
  wire n18933_o;
  reg n18934_q;
  wire n18935_o;
  wire n18936_o;
  reg n18937_q;
  wire n18938_o;
  wire n18939_o;
  reg n18940_q;
  wire n18941_o;
  wire n18942_o;
  reg n18943_q;
  wire n18944_o;
  wire n18945_o;
  reg n18946_q;
  wire n18947_o;
  wire n18948_o;
  reg n18949_q;
  wire n18950_o;
  wire n18951_o;
  reg n18952_q;
  wire n18953_o;
  wire n18954_o;
  reg n18955_q;
  wire [48:0] n18956_o;
  wire [5:0] nie_block_wl;
  wire [1:0] n18957_o;
  wire [2:0] n18958_o;
  wire [3:0] n18959_o;
  wire [4:0] n18960_o;
  wire [5:0] n18961_o;
  wire n18963_o;
  wire [2:0] n18965_o;
  wire n18966_o;
  wire [3:0] n18967_o;
  wire n18968_o;
  wire [4:0] n18969_o;
  wire n18970_o;
  wire [5:0] n18971_o;
  wire n18977_o;
  wire n18978_o;
  wire n18979_o;
  wire n18981_o;
  wire n18983_o;
  wire n18984_o;
  wire n18985_o;
  wire n18986_o;
  wire n18987_o;
  wire n18988_o;
  wire n18989_o;
  wire n18990_o;
  wire n18991_o;
  wire n18992_o;
  wire n18993_o;
  wire n18994_o;
  wire n18995_o;
  wire n18996_o;
  wire n18997_o;
  wire n18998_o;
  wire n18999_o;
  wire n19000_o;
  wire n19001_o;
  wire n19002_o;
  wire n19003_o;
  wire n19005_o;
  wire n19006_o;
  wire n19007_o;
  wire [1:0] n19008_o;
  wire n19009_o;
  wire [2:0] n19010_o;
  wire n19011_o;
  wire [3:0] n19012_o;
  wire n19013_o;
  wire [4:0] n19014_o;
  wire n19015_o;
  wire [5:0] n19016_o;
  wire n19022_o;
  wire n19023_o;
  wire n19024_o;
  wire n19026_o;
  wire n19028_o;
  wire n19029_o;
  wire n19030_o;
  wire n19031_o;
  wire n19032_o;
  wire n19033_o;
  wire n19034_o;
  wire n19035_o;
  wire n19036_o;
  wire n19037_o;
  wire n19038_o;
  wire n19039_o;
  wire n19040_o;
  wire n19041_o;
  wire n19042_o;
  wire n19043_o;
  wire n19044_o;
  wire n19045_o;
  wire n19046_o;
  wire n19047_o;
  wire n19048_o;
  wire n19050_o;
  wire n19051_o;
  wire n19052_o;
  wire [1:0] n19053_o;
  wire n19054_o;
  wire [2:0] n19055_o;
  wire n19056_o;
  wire [3:0] n19057_o;
  wire n19058_o;
  wire [4:0] n19059_o;
  wire n19060_o;
  wire [5:0] n19061_o;
  wire n19067_o;
  wire n19068_o;
  wire n19069_o;
  wire n19071_o;
  wire n19073_o;
  wire n19074_o;
  wire n19075_o;
  wire n19076_o;
  wire n19077_o;
  wire n19078_o;
  wire n19079_o;
  wire n19080_o;
  wire n19081_o;
  wire n19082_o;
  wire n19083_o;
  wire n19084_o;
  wire n19085_o;
  wire n19086_o;
  wire n19087_o;
  wire n19088_o;
  wire n19089_o;
  wire n19090_o;
  wire n19091_o;
  wire n19092_o;
  wire n19093_o;
  wire n19095_o;
  wire n19096_o;
  wire n19097_o;
  wire [1:0] n19098_o;
  wire n19099_o;
  wire [2:0] n19100_o;
  wire n19101_o;
  wire [3:0] n19102_o;
  wire n19103_o;
  wire [4:0] n19104_o;
  wire n19105_o;
  wire [5:0] n19106_o;
  wire n19112_o;
  wire n19113_o;
  wire n19114_o;
  wire n19116_o;
  wire n19118_o;
  wire n19119_o;
  wire n19120_o;
  wire n19121_o;
  wire n19122_o;
  wire n19123_o;
  wire n19124_o;
  wire n19125_o;
  wire n19126_o;
  wire n19127_o;
  wire n19128_o;
  wire n19129_o;
  wire n19130_o;
  wire n19131_o;
  wire n19132_o;
  wire n19133_o;
  wire n19134_o;
  wire n19135_o;
  wire n19136_o;
  wire n19137_o;
  wire n19138_o;
  wire n19140_o;
  wire n19141_o;
  wire n19142_o;
  wire [1:0] n19143_o;
  wire n19144_o;
  wire [2:0] n19145_o;
  wire n19146_o;
  wire [3:0] n19147_o;
  wire n19148_o;
  wire [4:0] n19149_o;
  wire n19150_o;
  wire [5:0] n19151_o;
  wire n19157_o;
  wire n19158_o;
  wire n19159_o;
  wire n19161_o;
  wire n19163_o;
  wire n19164_o;
  wire n19165_o;
  wire n19166_o;
  wire n19167_o;
  wire n19168_o;
  wire n19169_o;
  wire n19170_o;
  wire n19171_o;
  wire n19172_o;
  wire n19173_o;
  wire n19174_o;
  wire n19175_o;
  wire n19176_o;
  wire n19177_o;
  wire n19178_o;
  wire n19179_o;
  wire n19180_o;
  wire n19181_o;
  wire n19182_o;
  wire n19183_o;
  wire n19185_o;
  wire n19186_o;
  wire n19187_o;
  wire [1:0] n19188_o;
  wire n19189_o;
  wire [2:0] n19190_o;
  wire n19191_o;
  wire [3:0] n19192_o;
  wire n19193_o;
  wire [4:0] n19194_o;
  wire n19195_o;
  wire [5:0] n19196_o;
  wire n19202_o;
  wire n19203_o;
  wire n19204_o;
  wire n19206_o;
  wire n19208_o;
  wire n19209_o;
  wire n19210_o;
  wire n19211_o;
  wire n19212_o;
  wire n19213_o;
  wire n19214_o;
  wire n19215_o;
  wire n19216_o;
  wire n19217_o;
  wire n19218_o;
  wire n19219_o;
  wire n19220_o;
  wire n19221_o;
  wire n19222_o;
  wire n19223_o;
  wire n19224_o;
  wire n19225_o;
  wire n19226_o;
  wire n19227_o;
  wire n19228_o;
  wire n19230_o;
  wire n19231_o;
  wire n19232_o;
  wire [1:0] n19233_o;
  wire n19234_o;
  wire [2:0] n19235_o;
  wire n19236_o;
  wire [3:0] n19237_o;
  wire n19238_o;
  wire [4:0] n19239_o;
  wire n19240_o;
  wire [5:0] n19241_o;
  wire n19247_o;
  wire n19248_o;
  wire n19249_o;
  wire n19251_o;
  wire n19253_o;
  wire n19254_o;
  wire n19255_o;
  wire n19256_o;
  wire n19257_o;
  wire n19258_o;
  wire n19259_o;
  wire n19260_o;
  wire n19261_o;
  wire n19262_o;
  wire n19263_o;
  wire n19264_o;
  wire n19265_o;
  wire n19266_o;
  wire n19267_o;
  wire n19268_o;
  wire n19269_o;
  wire n19270_o;
  wire n19271_o;
  wire n19272_o;
  wire n19273_o;
  wire n19275_o;
  wire n19276_o;
  wire n19277_o;
  wire [1:0] n19278_o;
  wire n19279_o;
  wire [2:0] n19280_o;
  wire n19281_o;
  wire [3:0] n19282_o;
  wire n19283_o;
  wire [4:0] n19284_o;
  wire n19285_o;
  wire [5:0] n19286_o;
  wire n19292_o;
  wire n19293_o;
  wire n19294_o;
  wire n19296_o;
  wire n19298_o;
  wire n19299_o;
  wire n19300_o;
  wire n19301_o;
  wire n19302_o;
  wire n19303_o;
  wire n19304_o;
  wire n19305_o;
  wire n19306_o;
  wire n19307_o;
  wire n19308_o;
  wire n19309_o;
  wire n19310_o;
  wire n19311_o;
  wire n19312_o;
  wire n19313_o;
  wire n19314_o;
  wire n19315_o;
  wire n19316_o;
  wire n19317_o;
  wire n19318_o;
  wire n19320_o;
  wire n19321_o;
  wire n19322_o;
  wire [1:0] n19323_o;
  wire n19324_o;
  wire [2:0] n19325_o;
  wire n19326_o;
  wire [3:0] n19327_o;
  wire n19328_o;
  wire [4:0] n19329_o;
  wire n19330_o;
  wire [5:0] n19331_o;
  wire n19337_o;
  wire n19338_o;
  wire n19339_o;
  wire n19341_o;
  wire n19343_o;
  wire n19344_o;
  wire n19345_o;
  wire n19346_o;
  wire n19347_o;
  wire n19348_o;
  wire n19349_o;
  wire n19350_o;
  wire n19351_o;
  wire n19352_o;
  wire n19353_o;
  wire n19354_o;
  wire n19355_o;
  wire n19356_o;
  wire n19357_o;
  wire n19358_o;
  wire n19359_o;
  wire n19360_o;
  wire n19361_o;
  wire n19362_o;
  wire n19363_o;
  wire n19365_o;
  wire [2:0] n19367_o;
  wire n19368_o;
  wire [3:0] n19369_o;
  wire n19370_o;
  wire [4:0] n19371_o;
  wire n19372_o;
  wire [5:0] n19373_o;
  wire n19379_o;
  wire n19380_o;
  wire n19381_o;
  wire n19383_o;
  wire n19385_o;
  wire n19386_o;
  wire n19387_o;
  wire n19388_o;
  wire n19389_o;
  wire n19390_o;
  wire n19391_o;
  wire n19392_o;
  wire n19393_o;
  wire n19394_o;
  wire n19395_o;
  wire n19396_o;
  wire n19397_o;
  wire n19398_o;
  wire n19399_o;
  wire n19400_o;
  wire n19401_o;
  wire n19402_o;
  wire n19403_o;
  wire n19404_o;
  wire n19405_o;
  wire n19407_o;
  wire [2:0] n19409_o;
  wire n19410_o;
  wire [3:0] n19411_o;
  wire n19412_o;
  wire [4:0] n19413_o;
  wire n19414_o;
  wire [5:0] n19415_o;
  wire n19421_o;
  wire n19422_o;
  wire n19423_o;
  wire n19425_o;
  wire n19427_o;
  wire n19428_o;
  wire n19429_o;
  wire n19430_o;
  wire n19431_o;
  wire n19432_o;
  wire n19433_o;
  wire n19434_o;
  wire n19435_o;
  wire n19436_o;
  wire n19437_o;
  wire n19438_o;
  wire n19439_o;
  wire n19440_o;
  wire n19441_o;
  wire n19442_o;
  wire n19443_o;
  wire n19444_o;
  wire n19445_o;
  wire n19446_o;
  wire n19447_o;
  wire n19449_o;
  wire [2:0] n19451_o;
  wire n19452_o;
  wire [3:0] n19453_o;
  wire n19454_o;
  wire [4:0] n19455_o;
  wire n19456_o;
  wire [5:0] n19457_o;
  wire n19463_o;
  wire n19464_o;
  wire n19465_o;
  wire n19467_o;
  wire n19469_o;
  wire n19470_o;
  wire n19471_o;
  wire n19472_o;
  wire n19473_o;
  wire n19474_o;
  wire n19475_o;
  wire n19476_o;
  wire n19477_o;
  wire n19478_o;
  wire n19479_o;
  wire n19480_o;
  wire n19481_o;
  wire n19482_o;
  wire n19483_o;
  wire n19484_o;
  wire n19485_o;
  wire n19486_o;
  wire n19487_o;
  wire n19488_o;
  wire n19489_o;
  wire dac_block_pwmsel;
  wire dac_block_pwm_block_pwm0;
  wire dac_block_pwm_block_pwm1;
  wire dac_block_pwm_block_pwm2;
  wire dac_block_pwm_block_nc2d10xr9del;
  wire dac_block_pwm_block_pwmreg1toggle;
  wire dac_block_pwm_block_pwmreg2toggle;
  wire dac_block_pwm_block_pwmreg0;
  wire dac_block_pwm_block_pwmreg1;
  wire dac_block_pwm_block_pwmreg2;
  wire dac_block_pwm_block_pwmcomm;
  wire dac_block_pwm_block_pwmcommdel;
  wire dac_block_pwm_block_pwmcommand;
  wire dac_block_pwm_block_pwmcomp;
  wire n19490_o;
  wire n19491_o;
  wire n19492_o;
  wire n19493_o;
  wire n19494_o;
  wire n19495_o;
  wire n19496_o;
  wire n19497_o;
  wire n19498_o;
  wire n19499_o;
  wire n19500_o;
  wire n19501_o;
  wire dac_block_pwm_block_nc2d10xr9del_b_o_out;
  wire n19502_o;
  wire n19503_o;
  wire n19504_o;
  wire n19505_o;
  wire n19506_o;
  wire n19508_o;
  wire n19509_o;
  wire n19510_o;
  wire n19518_o;
  wire n19520_o;
  wire n19522_o;
  wire n19523_o;
  wire n19524_o;
  wire n19525_o;
  wire n19526_o;
  wire n19527_o;
  wire n19529_o;
  wire n19531_o;
  wire n19533_o;
  wire [1:0] n19539_o;
  wire [2:0] n19540_o;
  wire n19546_o;
  wire n19548_o;
  wire n19550_o;
  wire n19551_o;
  wire n19552_o;
  wire n19553_o;
  wire n19554_o;
  wire dac_block_pwm_block_pwmcommdel_b_o_out;
  wire n19555_o;
  wire n19556_o;
  wire n19557_o;
  wire n19558_o;
  wire n19560_o;
  wire [1:0] n19562_o;
  wire [2:0] n19563_o;
  wire [1:0] n19564_o;
  wire [2:0] n19565_o;
  wire n19571_o;
  wire n19572_o;
  wire n19573_o;
  wire n19574_o;
  wire n19576_o;
  wire n19578_o;
  wire n19579_o;
  wire n19580_o;
  wire n19581_o;
  wire n19582_o;
  wire n19583_o;
  wire n19584_o;
  wire n19585_o;
  wire n19586_o;
  wire n19587_o;
  wire n19588_o;
  wire dac_block_pwm_block_pwmsr_b_o_q;
  wire n19589_o;
  wire n19591_o;
  wire n19592_o;
  wire n19593_o;
  wire n19594_o;
  reg n19595_q;
  wire n19596_o;
  reg n19597_q;
  wire n19598_o;
  reg n19599_q;
  wire [4:0] dac_block_dacrom_block_ndac;
  wire [6:0] dac_block_dacrom_block_dacval;
  wire [6:0] dac_block_dacrom_block_dacpwm;
  wire n19600_o;
  wire [3:0] n19601_o;
  wire [3:0] n19602_o;
  wire [4:0] n19603_o;
  wire n19604_o;
  wire [4:0] n19605_o;
  wire n19606_o;
  wire [3:0] n19607_o;
  wire [3:0] n19608_o;
  wire [4:0] n19609_o;
  wire [4:0] n19610_o;
  wire [6:0] n19611_o;
  wire [6:0] n19613_o;
  wire [6:0] n19615_o;
  wire [6:0] n19616_o;
  wire [6:0] n19618_o;
  wire [5:0] n19619_o;
  localparam n19620_o = 1'b0;
  wire [5:0] abus_block_wl;
  wire [1:0] n19621_o;
  wire [2:0] n19622_o;
  wire [3:0] n19623_o;
  wire [4:0] n19624_o;
  wire [5:0] n19625_o;
  wire n19627_o;
  wire n19628_o;
  wire [1:0] n19629_o;
  wire n19630_o;
  wire n19631_o;
  wire [2:0] n19632_o;
  wire n19633_o;
  wire n19634_o;
  wire [3:0] n19635_o;
  wire [4:0] n19637_o;
  wire [5:0] n19639_o;
  wire n19645_o;
  wire n19646_o;
  wire n19647_o;
  wire n19649_o;
  wire n19651_o;
  wire n19652_o;
  wire n19653_o;
  wire n19654_o;
  wire n19655_o;
  wire n19656_o;
  wire n19657_o;
  wire n19658_o;
  wire n19659_o;
  wire n19660_o;
  wire n19661_o;
  wire n19662_o;
  wire n19663_o;
  wire n19664_o;
  wire n19665_o;
  wire n19666_o;
  wire n19667_o;
  wire n19668_o;
  wire n19669_o;
  wire n19670_o;
  wire n19671_o;
  wire n19672_o;
  wire n19674_o;
  wire n19675_o;
  wire [1:0] n19676_o;
  wire n19677_o;
  wire n19678_o;
  wire [2:0] n19679_o;
  wire n19680_o;
  wire n19681_o;
  wire [3:0] n19682_o;
  wire [4:0] n19684_o;
  wire [5:0] n19686_o;
  wire n19692_o;
  wire n19693_o;
  wire n19694_o;
  wire n19696_o;
  wire n19698_o;
  wire n19699_o;
  wire n19700_o;
  wire n19701_o;
  wire n19702_o;
  wire n19703_o;
  wire n19704_o;
  wire n19705_o;
  wire n19706_o;
  wire n19707_o;
  wire n19708_o;
  wire n19709_o;
  wire n19710_o;
  wire n19711_o;
  wire n19712_o;
  wire n19713_o;
  wire n19714_o;
  wire n19715_o;
  wire n19716_o;
  wire n19717_o;
  wire n19718_o;
  wire n19719_o;
  wire n19721_o;
  wire n19722_o;
  wire [1:0] n19723_o;
  wire n19724_o;
  wire n19725_o;
  wire [2:0] n19726_o;
  wire n19727_o;
  wire n19728_o;
  wire [3:0] n19729_o;
  wire [4:0] n19731_o;
  wire [5:0] n19733_o;
  wire n19739_o;
  wire n19740_o;
  wire n19741_o;
  wire n19743_o;
  wire n19745_o;
  wire n19746_o;
  wire n19747_o;
  wire n19748_o;
  wire n19749_o;
  wire n19750_o;
  wire n19751_o;
  wire n19752_o;
  wire n19753_o;
  wire n19754_o;
  wire n19755_o;
  wire n19756_o;
  wire n19757_o;
  wire n19758_o;
  wire n19759_o;
  wire n19760_o;
  wire n19761_o;
  wire n19762_o;
  wire n19763_o;
  wire n19764_o;
  wire n19765_o;
  wire n19766_o;
  wire n19768_o;
  wire n19769_o;
  wire [1:0] n19770_o;
  wire n19771_o;
  wire n19772_o;
  wire [2:0] n19773_o;
  wire n19774_o;
  wire n19775_o;
  wire [3:0] n19776_o;
  wire [4:0] n19778_o;
  wire [5:0] n19780_o;
  wire n19786_o;
  wire n19787_o;
  wire n19788_o;
  wire n19790_o;
  wire n19792_o;
  wire n19793_o;
  wire n19794_o;
  wire n19795_o;
  wire n19796_o;
  wire n19797_o;
  wire n19798_o;
  wire n19799_o;
  wire n19800_o;
  wire n19801_o;
  wire n19802_o;
  wire n19803_o;
  wire n19804_o;
  wire n19805_o;
  wire n19806_o;
  wire n19807_o;
  wire n19808_o;
  wire n19809_o;
  wire n19810_o;
  wire n19811_o;
  wire n19812_o;
  wire n19813_o;
  wire n19815_o;
  wire n19816_o;
  wire [1:0] n19817_o;
  wire n19818_o;
  wire n19819_o;
  wire [2:0] n19820_o;
  wire n19821_o;
  wire n19822_o;
  wire [3:0] n19823_o;
  wire [4:0] n19825_o;
  wire [5:0] n19827_o;
  wire n19833_o;
  wire n19834_o;
  wire n19835_o;
  wire n19837_o;
  wire n19839_o;
  wire n19840_o;
  wire n19841_o;
  wire n19842_o;
  wire n19843_o;
  wire n19844_o;
  wire n19845_o;
  wire n19846_o;
  wire n19847_o;
  wire n19848_o;
  wire n19849_o;
  wire n19850_o;
  wire n19851_o;
  wire n19852_o;
  wire n19853_o;
  wire n19854_o;
  wire n19855_o;
  wire n19856_o;
  wire n19857_o;
  wire n19858_o;
  wire n19859_o;
  wire n19860_o;
  wire n19862_o;
  wire n19863_o;
  wire [1:0] n19864_o;
  wire n19865_o;
  wire n19866_o;
  wire [2:0] n19867_o;
  wire n19868_o;
  wire n19869_o;
  wire [3:0] n19870_o;
  wire [4:0] n19872_o;
  wire [5:0] n19874_o;
  wire n19880_o;
  wire n19881_o;
  wire n19882_o;
  wire n19884_o;
  wire n19886_o;
  wire n19887_o;
  wire n19888_o;
  wire n19889_o;
  wire n19890_o;
  wire n19891_o;
  wire n19892_o;
  wire n19893_o;
  wire n19894_o;
  wire n19895_o;
  wire n19896_o;
  wire n19897_o;
  wire n19898_o;
  wire n19899_o;
  wire n19900_o;
  wire n19901_o;
  wire n19902_o;
  wire n19903_o;
  wire n19904_o;
  wire n19905_o;
  wire n19906_o;
  wire n19907_o;
  wire n19909_o;
  wire n19910_o;
  wire [1:0] n19911_o;
  wire n19912_o;
  wire n19913_o;
  wire [2:0] n19914_o;
  wire n19915_o;
  wire n19916_o;
  wire [3:0] n19917_o;
  wire [4:0] n19919_o;
  wire [5:0] n19921_o;
  wire n19927_o;
  wire n19928_o;
  wire n19929_o;
  wire n19931_o;
  wire n19933_o;
  wire n19934_o;
  wire n19935_o;
  wire n19936_o;
  wire n19937_o;
  wire n19938_o;
  wire n19939_o;
  wire n19940_o;
  wire n19941_o;
  wire n19942_o;
  wire n19943_o;
  wire n19944_o;
  wire n19945_o;
  wire n19946_o;
  wire n19947_o;
  wire n19948_o;
  wire n19949_o;
  wire n19950_o;
  wire n19951_o;
  wire n19952_o;
  wire n19953_o;
  wire n19954_o;
  wire n19956_o;
  wire n19957_o;
  wire [1:0] n19958_o;
  wire n19959_o;
  wire n19960_o;
  wire [2:0] n19961_o;
  wire n19962_o;
  wire n19963_o;
  wire [3:0] n19964_o;
  wire [4:0] n19966_o;
  wire [5:0] n19968_o;
  wire n19974_o;
  wire n19975_o;
  wire n19976_o;
  wire n19978_o;
  wire n19980_o;
  wire n19981_o;
  wire n19982_o;
  wire n19983_o;
  wire n19984_o;
  wire n19985_o;
  wire n19986_o;
  wire n19987_o;
  wire n19988_o;
  wire n19989_o;
  wire n19990_o;
  wire n19991_o;
  wire n19992_o;
  wire n19993_o;
  wire n19994_o;
  wire n19995_o;
  wire n19996_o;
  wire n19997_o;
  wire n19998_o;
  wire n19999_o;
  wire n20000_o;
  wire n20001_o;
  wire n20003_o;
  wire n20004_o;
  wire [1:0] n20005_o;
  wire n20006_o;
  wire n20007_o;
  wire [2:0] n20008_o;
  wire n20009_o;
  wire n20010_o;
  wire [3:0] n20011_o;
  wire [4:0] n20013_o;
  wire [5:0] n20015_o;
  wire n20021_o;
  wire n20022_o;
  wire n20023_o;
  wire n20025_o;
  wire n20027_o;
  wire n20028_o;
  wire n20029_o;
  wire n20030_o;
  wire n20031_o;
  wire n20032_o;
  wire n20033_o;
  wire n20034_o;
  wire n20035_o;
  wire n20036_o;
  wire n20037_o;
  wire n20038_o;
  wire n20039_o;
  wire n20040_o;
  wire n20041_o;
  wire n20042_o;
  wire n20043_o;
  wire n20044_o;
  wire n20045_o;
  wire n20046_o;
  wire n20047_o;
  wire n20048_o;
  wire n20050_o;
  wire n20051_o;
  wire n20052_o;
  wire [1:0] n20053_o;
  wire n20054_o;
  wire n20055_o;
  wire [2:0] n20056_o;
  wire n20057_o;
  wire n20058_o;
  wire [3:0] n20059_o;
  wire [4:0] n20061_o;
  wire [5:0] n20063_o;
  wire n20069_o;
  wire n20070_o;
  wire n20071_o;
  wire n20073_o;
  wire n20075_o;
  wire n20076_o;
  wire n20077_o;
  wire n20078_o;
  wire n20079_o;
  wire n20080_o;
  wire n20081_o;
  wire n20082_o;
  wire n20083_o;
  wire n20084_o;
  wire n20085_o;
  wire n20086_o;
  wire n20087_o;
  wire n20088_o;
  wire n20089_o;
  wire n20090_o;
  wire n20091_o;
  wire n20092_o;
  wire n20093_o;
  wire n20094_o;
  wire n20095_o;
  wire n20096_o;
  wire n20098_o;
  wire [1:0] n20099_o;
  wire [2:0] n20101_o;
  wire [3:0] n20103_o;
  wire n20104_o;
  wire [4:0] n20105_o;
  wire [5:0] n20106_o;
  wire n20112_o;
  wire n20113_o;
  wire n20114_o;
  wire n20116_o;
  wire n20118_o;
  wire n20119_o;
  wire n20120_o;
  wire n20121_o;
  wire n20122_o;
  wire n20123_o;
  wire n20124_o;
  wire n20125_o;
  wire n20126_o;
  wire n20127_o;
  wire n20128_o;
  wire n20129_o;
  wire n20130_o;
  wire n20131_o;
  wire n20132_o;
  wire n20133_o;
  wire n20134_o;
  wire n20135_o;
  wire n20136_o;
  wire n20137_o;
  wire n20138_o;
  wire n20139_o;
  wire n20141_o;
  wire [1:0] n20142_o;
  wire [2:0] n20144_o;
  wire [3:0] n20146_o;
  wire [4:0] n20147_o;
  wire [5:0] n20149_o;
  wire n20155_o;
  wire n20156_o;
  wire n20157_o;
  wire n20159_o;
  wire n20161_o;
  wire n20162_o;
  wire n20163_o;
  wire n20164_o;
  wire n20165_o;
  wire n20166_o;
  wire n20167_o;
  wire n20168_o;
  wire n20169_o;
  wire n20170_o;
  wire n20171_o;
  wire n20172_o;
  wire n20173_o;
  wire n20174_o;
  wire n20175_o;
  wire n20176_o;
  wire n20177_o;
  wire n20178_o;
  wire n20179_o;
  wire n20180_o;
  wire n20181_o;
  wire n20182_o;
  wire n20184_o;
  wire n20185_o;
  wire [1:0] n20186_o;
  wire [2:0] n20188_o;
  wire n20189_o;
  wire n20190_o;
  wire [3:0] n20191_o;
  wire n20192_o;
  wire [4:0] n20193_o;
  wire [5:0] n20195_o;
  wire n20201_o;
  wire n20202_o;
  wire n20203_o;
  wire n20205_o;
  wire n20207_o;
  wire n20208_o;
  wire n20209_o;
  wire n20210_o;
  wire n20211_o;
  wire n20212_o;
  wire n20213_o;
  wire n20214_o;
  wire n20215_o;
  wire n20216_o;
  wire n20217_o;
  wire n20218_o;
  wire n20219_o;
  wire n20220_o;
  wire n20221_o;
  wire n20222_o;
  wire n20223_o;
  wire n20224_o;
  wire n20225_o;
  wire n20226_o;
  wire n20227_o;
  wire n20228_o;
  wire n20230_o;
  wire n20231_o;
  wire [1:0] n20232_o;
  wire [2:0] n20234_o;
  wire n20235_o;
  wire n20236_o;
  wire [3:0] n20237_o;
  wire [4:0] n20238_o;
  wire [5:0] n20240_o;
  wire n20246_o;
  wire n20247_o;
  wire n20248_o;
  wire n20250_o;
  wire n20252_o;
  wire n20253_o;
  wire n20254_o;
  wire n20255_o;
  wire n20256_o;
  wire n20257_o;
  wire n20258_o;
  wire n20259_o;
  wire n20260_o;
  wire n20261_o;
  wire n20262_o;
  wire n20263_o;
  wire n20264_o;
  wire n20265_o;
  wire n20266_o;
  wire n20267_o;
  wire n20268_o;
  wire n20269_o;
  wire n20270_o;
  wire n20271_o;
  wire n20272_o;
  wire n20273_o;
  wire n20275_o;
  wire [1:0] n20277_o;
  wire [2:0] n20279_o;
  wire [3:0] n20281_o;
  wire [4:0] n20282_o;
  wire [5:0] n20284_o;
  wire n20290_o;
  wire n20291_o;
  wire n20292_o;
  wire n20294_o;
  wire n20296_o;
  wire n20297_o;
  wire n20298_o;
  wire n20299_o;
  wire n20300_o;
  wire n20301_o;
  wire n20302_o;
  wire n20303_o;
  wire n20304_o;
  wire n20305_o;
  wire n20306_o;
  wire n20307_o;
  wire n20308_o;
  wire n20309_o;
  wire n20310_o;
  wire n20311_o;
  wire n20312_o;
  wire n20313_o;
  wire n20314_o;
  wire n20315_o;
  wire n20316_o;
  wire n20317_o;
  wire n20319_o;
  wire [1:0] n20321_o;
  wire [2:0] n20323_o;
  wire [3:0] n20325_o;
  wire [4:0] n20327_o;
  wire [5:0] n20329_o;
  wire n20335_o;
  wire n20336_o;
  wire n20337_o;
  wire n20339_o;
  wire n20341_o;
  wire n20342_o;
  wire n20343_o;
  wire n20344_o;
  wire n20345_o;
  wire n20346_o;
  wire n20347_o;
  wire n20348_o;
  wire n20349_o;
  wire n20350_o;
  wire n20351_o;
  wire n20352_o;
  wire n20353_o;
  wire n20354_o;
  wire n20355_o;
  wire n20356_o;
  wire n20357_o;
  wire n20358_o;
  wire n20359_o;
  wire n20360_o;
  wire n20361_o;
  wire n20362_o;
  wire [9:0] n20363_o;
  wire n20364_o;
  wire [9:0] n20365_o;
  wire [9:0] n20366_o;
  wire [9:0] n20367_o;
  wire n20368_o;
  wire n20369_o;
  wire mte_delay_b_o_out;
  wire n20370_o;
  wire n20371_o;
  wire n20372_o;
  wire n20373_o;
  wire n20374_o;
  wire n20376_o;
  wire n20377_o;
  wire n20378_o;
  reg n20379_q;
  wire [3:0] n20380_o;
  wire [7:0] n20381_o;
  wire [10:0] n20382_o;
  reg [10:0] n20383_q;
  wire n20384_o;
  reg n20385_q;
  wire [7:0] n20386_o;
  reg [7:0] n20387_q;
  wire [15:0] n20388_o;
  reg [15:0] n20389_q;
  wire [4:0] n20390_o;
  wire [9:0] n20391_o;
  wire [11:0] n20392_o;
  wire [7:0] n20393_o;
  reg [7:0] n20394_q;
  wire [11:0] n20395_o;
  wire [11:0] n20396_o;
  reg [11:0] n20397_q;
  wire [15:0] n20398_o;
  wire [9:0] n20400_data; // mem_rd
  wire [11:0] n20403_data; // mem_rd
  wire [11:0] n20406_data; // mem_rd
  wire n20408_o;
  wire n20409_o;
  wire n20410_o;
  wire n20411_o;
  wire n20412_o;
  wire n20413_o;
  wire n20414_o;
  wire n20415_o;
  wire n20416_o;
  wire n20417_o;
  wire n20418_o;
  wire n20419_o;
  wire n20420_o;
  wire n20421_o;
  wire n20422_o;
  wire n20423_o;
  wire n20424_o;
  wire n20425_o;
  wire n20426_o;
  wire n20427_o;
  wire n20428_o;
  wire n20429_o;
  wire n20430_o;
  wire n20431_o;
  wire n20432_o;
  wire n20433_o;
  wire n20434_o;
  wire n20435_o;
  wire n20436_o;
  wire n20437_o;
  wire n20438_o;
  wire n20439_o;
  wire n20440_o;
  wire n20441_o;
  wire n20442_o;
  wire n20443_o;
  wire n20444_o;
  wire n20445_o;
  wire n20446_o;
  wire n20447_o;
  wire n20448_o;
  wire n20449_o;
  wire n20450_o;
  wire n20451_o;
  wire n20452_o;
  wire n20453_o;
  wire n20454_o;
  wire n20455_o;
  wire n20456_o;
  wire n20457_o;
  wire n20458_o;
  wire n20459_o;
  wire n20460_o;
  wire n20461_o;
  wire n20462_o;
  wire n20463_o;
  wire n20464_o;
  wire n20465_o;
  wire n20466_o;
  wire n20467_o;
  wire n20468_o;
  wire n20469_o;
  wire n20470_o;
  wire n20471_o;
  wire n20472_o;
  wire n20473_o;
  wire n20474_o;
  wire n20475_o;
  wire n20476_o;
  wire n20477_o;
  wire n20478_o;
  wire n20479_o;
  wire n20480_o;
  wire n20481_o;
  wire n20482_o;
  wire n20483_o;
  wire n20484_o;
  wire n20485_o;
  wire n20486_o;
  wire n20487_o;
  wire n20488_o;
  wire n20489_o;
  wire n20490_o;
  wire n20491_o;
  wire n20492_o;
  wire n20493_o;
  wire n20494_o;
  wire n20495_o;
  wire n20496_o;
  wire n20497_o;
  wire n20498_o;
  wire n20499_o;
  wire n20500_o;
  wire n20501_o;
  wire n20502_o;
  wire n20503_o;
  wire n20504_o;
  wire n20505_o;
  wire n20506_o;
  wire n20507_o;
  wire n20508_o;
  wire n20509_o;
  wire n20510_o;
  wire n20511_o;
  wire n20512_o;
  wire n20513_o;
  wire n20514_o;
  wire n20515_o;
  wire n20516_o;
  wire n20517_o;
  wire n20518_o;
  wire n20519_o;
  wire n20520_o;
  wire n20521_o;
  wire n20522_o;
  wire n20523_o;
  wire n20524_o;
  wire n20525_o;
  wire n20526_o;
  wire n20527_o;
  wire n20528_o;
  wire n20529_o;
  wire n20530_o;
  wire n20531_o;
  wire n20532_o;
  wire n20533_o;
  wire n20534_o;
  wire n20535_o;
  wire n20536_o;
  wire n20537_o;
  wire n20538_o;
  wire n20539_o;
  wire n20540_o;
  wire n20541_o;
  wire [31:0] n20542_o;
  wire n20543_o;
  wire n20544_o;
  wire n20545_o;
  wire n20546_o;
  wire n20547_o;
  wire n20548_o;
  wire n20549_o;
  wire n20550_o;
  wire n20551_o;
  wire n20552_o;
  wire n20553_o;
  wire n20554_o;
  wire n20555_o;
  wire n20556_o;
  wire n20557_o;
  wire n20558_o;
  wire n20559_o;
  wire n20560_o;
  wire n20561_o;
  wire n20562_o;
  wire n20563_o;
  wire n20564_o;
  wire n20565_o;
  wire n20566_o;
  wire n20567_o;
  wire n20568_o;
  wire n20569_o;
  wire n20570_o;
  wire n20571_o;
  wire n20572_o;
  wire n20573_o;
  wire n20574_o;
  wire n20575_o;
  wire n20576_o;
  wire n20577_o;
  wire n20578_o;
  wire n20579_o;
  wire n20580_o;
  wire n20581_o;
  wire n20582_o;
  wire n20583_o;
  wire n20584_o;
  wire n20585_o;
  wire n20586_o;
  wire n20587_o;
  wire n20588_o;
  wire n20589_o;
  wire n20590_o;
  wire n20591_o;
  wire n20592_o;
  wire n20593_o;
  wire n20594_o;
  wire n20595_o;
  wire [11:0] n20596_o;
  assign o_tst2 = n19620_o;
  assign o_tst4 = n119_o;
  assign o_a = n20398_o;
  assign o_me_l = n20369_o;
  assign o_mte = mte_delay_b_o_out;
  assign o_bsy = n20368_o;
  assign o_dao = n19619_o;
  assign o_audio = n20365_o;
  /* vlm5030_gl.vhd:164:10  */
  assign osc = n14_o; // (signal)
  /* vlm5030_gl.vhd:165:10  */
  always @*
    clk2 = n20380_o; // (isignal)
  initial
    clk2 = 4'b0000;
  /* vlm5030_gl.vhd:166:10  */
  assign nclk2 = n295_o; // (signal)
  /* vlm5030_gl.vhd:168:10  */
  assign rst = n123_o; // (signal)
  /* vlm5030_gl.vhd:171:10  */
  assign dq = n20381_o; // (signal)
  /* vlm5030_gl.vhd:172:10  */
  assign maskdq53 = dq_block_maskdq53s; // (signal)
  /* vlm5030_gl.vhd:174:10  */
  assign starttst = n217_o; // (signal)
  /* vlm5030_gl.vhd:175:10  */
  assign tststopclk2 = n222_o; // (signal)
  /* vlm5030_gl.vhd:175:23  */
  assign tstend2id = n225_o; // (signal)
  /* vlm5030_gl.vhd:175:34  */
  assign tstend2ie = n229_o; // (signal)
  /* vlm5030_gl.vhd:176:10  */
  assign tstenid2a = n232_o; // (signal)
  /* vlm5030_gl.vhd:176:21  */
  assign tstenie2a = n235_o; // (signal)
  /* vlm5030_gl.vhd:176:32  */
  assign tstenctrl2a = n239_o; // (signal)
  /* vlm5030_gl.vhd:177:10  */
  assign tstenie2dac = n242_o; // (signal)
  /* vlm5030_gl.vhd:179:10  */
  always @*
    clk2divq = n20383_q; // (isignal)
  initial
    clk2divq = 11'b00000000000;
  /* vlm5030_gl.vhd:180:10  */
  assign c2d0 = n358_o; // (signal)
  /* vlm5030_gl.vhd:180:16  */
  assign c2d1 = n375_o; // (signal)
  /* vlm5030_gl.vhd:181:10  */
  assign c2d3 = n392_o; // (signal)
  /* vlm5030_gl.vhd:181:16  */
  assign c2d4 = n409_o; // (signal)
  /* vlm5030_gl.vhd:181:22  */
  assign c2d5 = n426_o; // (signal)
  /* vlm5030_gl.vhd:182:10  */
  assign c2d6 = n443_o; // (signal)
  /* vlm5030_gl.vhd:182:16  */
  assign c2d7 = n460_o; // (signal)
  /* vlm5030_gl.vhd:182:22  */
  assign c2d8 = n477_o; // (signal)
  /* vlm5030_gl.vhd:183:10  */
  assign c2d9 = n494_o; // (signal)
  /* vlm5030_gl.vhd:183:16  */
  assign c2d10 = n511_o; // (signal)
  /* vlm5030_gl.vhd:184:10  */
  assign c2d5fin = n524_o; // (signal)
  /* vlm5030_gl.vhd:185:10  */
  assign c2d7fin = n538_o; // (signal)
  /* vlm5030_gl.vhd:185:19  */
  assign nc2d7fin = n550_o; // (signal)
  /* vlm5030_gl.vhd:186:10  */
  assign c2d9fin = n563_o; // (signal)
  /* vlm5030_gl.vhd:186:19  */
  assign nc2d9fin = n575_o; // (signal)
  /* vlm5030_gl.vhd:187:10  */
  assign clk2gd5 = n639_o; // (signal)
  /* vlm5030_gl.vhd:188:10  */
  assign nc2d1 = n650_o; // (signal)
  /* vlm5030_gl.vhd:188:17  */
  assign nc2d6 = n687_o; // (signal)
  /* vlm5030_gl.vhd:189:10  */
  assign nc2d8 = n698_o; // (signal)
  /* vlm5030_gl.vhd:189:17  */
  assign nc2d10 = n709_o; // (signal)
  /* vlm5030_gl.vhd:190:10  */
  assign c2d3gated = n676_o; // (signal)
  /* vlm5030_gl.vhd:193:10  */
  assign fsromevalout = n775_o; // (signal)
  /* vlm5030_gl.vhd:194:10  */
  assign fsromdo = n1952_o; // (signal)
  /* vlm5030_gl.vhd:195:10  */
  assign fsromnorhigh = n1974_o; // (signal)
  /* vlm5030_gl.vhd:196:10  */
  assign fsromnorlow = n1996_o; // (signal)
  /* vlm5030_gl.vhd:198:10  */
  assign clk2ctrl = n2021_o; // (signal)
  /* vlm5030_gl.vhd:199:10  */
  assign ncen1 = n2006_o; // (signal)
  /* vlm5030_gl.vhd:199:17  */
  assign cen3 = n2024_o; // (signal)
  /* vlm5030_gl.vhd:200:10  */
  assign eaoen = n2068_o; // (signal)
  /* vlm5030_gl.vhd:201:10  */
  always @*
    xromdo7nq = n20385_q; // (isignal)
  initial
    xromdo7nq = 1'b0;
  /* vlm5030_gl.vhd:202:10  */
  assign xromdo7q = n2063_o; // (signal)
  /* vlm5030_gl.vhd:203:10  */
  assign xromdo = n4216_o; // (signal)
  /* vlm5030_gl.vhd:204:10  */
  assign yromdo = n5046_o; // (signal)
  /* vlm5030_gl.vhd:205:10  */
  assign c2d3gate = n5045_o; // (signal)
  /* vlm5030_gl.vhd:208:10  */
  assign cntdn0 = n5074_o; // (signal)
  /* vlm5030_gl.vhd:211:10  */
  always @*
    dinalq = n20387_q; // (isignal)
  initial
    dinalq = 8'b00000000;
  /* vlm5030_gl.vhd:212:10  */
  assign aq = n20389_q; // (signal)
  /* vlm5030_gl.vhd:215:10  */
  assign startrise = n5260_o; // (signal)
  /* vlm5030_gl.vhd:216:10  */
  assign clkcntdn = n5622_o; // (signal)
  /* vlm5030_gl.vhd:217:10  */
  assign ncntdnload = n5560_o; // (signal)
  /* vlm5030_gl.vhd:218:10  */
  assign ncntdn = n5558_o; // (signal)
  /* vlm5030_gl.vhd:220:10  */
  assign eavcu = n5349_o; // (signal)
  /* vlm5030_gl.vhd:221:10  */
  assign ealatchh = n5368_o; // (signal)
  /* vlm5030_gl.vhd:222:10  */
  assign neaload = n5355_o; // (signal)
  /* vlm5030_gl.vhd:223:10  */
  assign eainc = n5630_o; // (signal)
  /* vlm5030_gl.vhd:224:10  */
  assign clrdinal = n5629_o; // (signal)
  /* vlm5030_gl.vhd:225:10  */
  assign clkdin = n5364_o; // (signal)
  /* vlm5030_gl.vhd:226:10  */
  assign nvcufinal = n5347_o; // (signal)
  /* vlm5030_gl.vhd:227:10  */
  assign vcufinal12 = n5343_o; // (signal)
  /* vlm5030_gl.vhd:228:10  */
  assign nbsy = n5669_o; // (signal)
  /* vlm5030_gl.vhd:229:10  */
  assign me = n5672_o; // (signal)
  /* vlm5030_gl.vhd:230:10  */
  assign rflatchwen = n5681_o; // (signal)
  /* vlm5030_gl.vhd:231:10  */
  assign asshift2 = n5686_o; // (signal)
  /* vlm5030_gl.vhd:232:10  */
  assign updtpitch = n5693_o; // (signal)
  /* vlm5030_gl.vhd:233:10  */
  assign enrf2id = n5703_o; // (signal)
  /* vlm5030_gl.vhd:234:10  */
  assign clkksa = start_block_n012x; // (signal)
  /* vlm5030_gl.vhd:235:10  */
  assign ensum2id = n5720_o; // (signal)
  /* vlm5030_gl.vhd:238:10  */
  assign clk2ena = n45_o; // (signal)
  /* vlm5030_gl.vhd:238:19  */
  assign clk2enb = n93_o; // (signal)
  /* vlm5030_gl.vhd:240:10  */
  assign rstdel = n138_o; // (signal)
  /* vlm5030_gl.vhd:243:10  */
  assign ksa = n20390_o; // (signal)
  /* vlm5030_gl.vhd:244:10  */
  assign nkdo = n12692_o; // (signal)
  /* vlm5030_gl.vhd:247:10  */
  assign rfdo = n13719_o; // (signal)
  /* vlm5030_gl.vhd:248:10  */
  assign rfdo97zero = n13735_o; // (signal)
  /* vlm5030_gl.vhd:251:10  */
  assign nid = n20391_o; // (signal)
  /* vlm5030_gl.vhd:253:10  */
  assign assum = n14424_o; // (signal)
  /* vlm5030_gl.vhd:255:10  */
  assign nie = n20392_o; // (signal)
  /* vlm5030_gl.vhd:257:10  */
  assign idlat = n20394_q; // (signal)
  /* vlm5030_gl.vhd:258:10  */
  assign idlatall1 = n15169_o; // (signal)
  /* vlm5030_gl.vhd:259:10  */
  assign enidlinv2id = n15116_o; // (signal)
  /* vlm5030_gl.vhd:260:10  */
  assign enidl2ie = n15135_o; // (signal)
  /* vlm5030_gl.vhd:261:10  */
  assign enidlinv2ie = n15130_o; // (signal)
  /* vlm5030_gl.vhd:264:10  */
  assign pitchoverflow = n14622_o; // (signal)
  /* vlm5030_gl.vhd:265:10  */
  assign enpitchlat = n14519_o; // (signal)
  /* vlm5030_gl.vhd:268:10  */
  assign enmem02id = n15203_o; // (signal)
  /* vlm5030_gl.vhd:269:10  */
  assign nmem0do = n15228_o; // (signal)
  /* vlm5030_gl.vhd:270:10  */
  assign mem0do = n15230_o; // (signal)
  /* vlm5030_gl.vhd:271:10  */
  assign enmem12ie = n15248_o; // (signal)
  /* vlm5030_gl.vhd:272:10  */
  assign mem1do2ie = n15273_o; // (signal)
  /* vlm5030_gl.vhd:273:10  */
  assign enmem22ie = n15293_o; // (signal)
  /* vlm5030_gl.vhd:274:10  */
  assign mem2do2ie = n15318_o; // (signal)
  /* vlm5030_gl.vhd:276:10  */
  assign ieregdrv = n18739_o; // (signal)
  /* vlm5030_gl.vhd:277:10  */
  assign ieregdrv4ie = n20395_o; // (signal)
  /* vlm5030_gl.vhd:278:10  */
  assign ieregload = n18867_o; // (signal)
  /* vlm5030_gl.vhd:280:10  */
  assign enieregfa2ie = n18877_o; // (signal)
  /* vlm5030_gl.vhd:282:10  */
  assign c2d10xr9 = n18891_o; // (signal)
  /* vlm5030_gl.vhd:283:10  */
  assign enie2a = n18892_o; // (signal)
  /* vlm5030_gl.vhd:284:10  */
  assign ieaddrreg = n20397_q; // (signal)
  /* vlm5030_gl.vhd:286:10  */
  assign pitchmod = n14640_o; // (signal)
  /* vlm5030_gl.vhd:288:10  */
  assign random = n5222_o; // (signal)
  /* vlm5030_gl.vhd:290:10  */
  assign pwmsr = dac_block_pwm_block_pwmsr_b_o_q; // (signal)
  assign n14_o = {1'b0, i_oscen, i_clk, i_clk};
  /* vlm5030_gl.vhd:304:28  */
  assign n17_o = ~(cen3 | tstenctrl2a);
  /* clock_functions_pack.vhd:139:26  */
  assign n22_o = clk2[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n23_o = clk2[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n24_o = n23_o | n17_o;
  /* clock_functions_pack.vhd:141:26  */
  assign n25_o = clk2[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n26_o = ~n17_o;
  /* clock_functions_pack.vhd:141:31  */
  assign n27_o = n25_o & n26_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n28_o = clk2[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n29_o = ~n17_o;
  /* clock_functions_pack.vhd:142:31  */
  assign n30_o = n28_o & n29_o;
  assign n31_o = {n30_o, n27_o, n24_o, n22_o};
  /* clock_functions_pack.vhd:139:26  */
  assign n36_o = n31_o[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n37_o = n31_o[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n38_o = n37_o | ncen1;
  /* clock_functions_pack.vhd:141:26  */
  assign n39_o = n31_o[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n40_o = ~ncen1;
  /* clock_functions_pack.vhd:141:31  */
  assign n41_o = n39_o & n40_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n42_o = n31_o[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n43_o = ~ncen1;
  /* clock_functions_pack.vhd:142:31  */
  assign n44_o = n42_o & n43_o;
  assign n45_o = {n44_o, n41_o, n38_o, n36_o};
  /* vlm5030_gl.vhd:305:28  */
  assign n49_o = ~(cen3 | tstenctrl2a);
  /* clock_functions_pack.vhd:139:26  */
  assign n54_o = clk2[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n55_o = clk2[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n56_o = n55_o | n49_o;
  /* clock_functions_pack.vhd:141:26  */
  assign n57_o = clk2[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n58_o = ~n49_o;
  /* clock_functions_pack.vhd:141:31  */
  assign n59_o = n57_o & n58_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n60_o = clk2[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n61_o = ~n49_o;
  /* clock_functions_pack.vhd:142:31  */
  assign n62_o = n60_o & n61_o;
  assign n63_o = {n62_o, n59_o, n56_o, n54_o};
  /* clock_functions_pack.vhd:139:26  */
  assign n68_o = n63_o[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n69_o = n63_o[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n70_o = n69_o | ncen1;
  /* clock_functions_pack.vhd:141:26  */
  assign n71_o = n63_o[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n72_o = ~ncen1;
  /* clock_functions_pack.vhd:141:31  */
  assign n73_o = n71_o & n72_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n74_o = n63_o[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n75_o = ~ncen1;
  /* clock_functions_pack.vhd:142:31  */
  assign n76_o = n74_o & n75_o;
  assign n77_o = {n76_o, n73_o, n70_o, n68_o};
  /* vlm5030_gl.vhd:305:65  */
  assign n78_o = fsromdo[6];
  /* vlm5030_gl.vhd:305:69  */
  assign n79_o = ~(n78_o | tstenctrl2a);
  /* clock_functions_pack.vhd:139:26  */
  assign n84_o = n77_o[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n85_o = n77_o[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n86_o = n85_o | n79_o;
  /* clock_functions_pack.vhd:141:26  */
  assign n87_o = n77_o[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n88_o = ~n79_o;
  /* clock_functions_pack.vhd:141:31  */
  assign n89_o = n87_o & n88_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n90_o = n77_o[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n91_o = ~n79_o;
  /* clock_functions_pack.vhd:142:31  */
  assign n92_o = n90_o & n91_o;
  assign n93_o = {n92_o, n89_o, n86_o, n84_o};
  /* vlm5030_gl.vhd:313:12  */
  always @*
    rstdel_block_porcnt = n141_q; // (isignal)
  initial
    rstdel_block_porcnt = 8'b11111111;
  /* vlm5030_gl.vhd:314:12  */
  always @*
    rstdel_block_npor = n143_q; // (isignal)
  initial
    rstdel_block_npor = 1'b0;
  /* vlm5030_gl.vhd:315:12  */
  always @*
    rstdel_block_del = n145_q; // (isignal)
  initial
    rstdel_block_del = 2'b00;
  assign n103_o = osc[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n105_o = osc[2];
  /* clock_functions_pack.vhd:65:34  */
  assign n106_o = n105_o & n113_o;
  /* vlm5030_gl.vhd:320:19  */
  assign n108_o = $unsigned(rstdel_block_porcnt) > $unsigned(8'b00000000);
  /* vlm5030_gl.vhd:321:28  */
  assign n110_o = rstdel_block_porcnt - 8'b00000001;
  /* vlm5030_gl.vhd:323:19  */
  assign n113_o = rstdel_block_porcnt == 8'b00000000;
  /* vlm5030_gl.vhd:329:15  */
  assign n119_o = ~rstdel_block_npor;
  /* vlm5030_gl.vhd:331:26  */
  assign n121_o = ~rstdel_block_npor;
  /* vlm5030_gl.vhd:331:32  */
  assign n122_o = n121_o & i_tst3;
  /* vlm5030_gl.vhd:331:16  */
  assign n123_o = n122_o ? 1'b1 : i_rst;
  assign n130_o = clk2[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n132_o = clk2[2];
  /* vlm5030_gl.vhd:336:19  */
  assign n134_o = rstdel_block_del[0];
  /* vlm5030_gl.vhd:336:23  */
  assign n135_o = {n134_o, rst};
  /* vlm5030_gl.vhd:340:18  */
  assign n138_o = rstdel_block_del[1];
  /* vlm5030_gl.vhd:319:7  */
  assign n139_o = n105_o & n108_o;
  /* vlm5030_gl.vhd:319:7  */
  assign n140_o = n139_o ? n110_o : rstdel_block_porcnt;
  /* vlm5030_gl.vhd:319:7  */
  always @(posedge n103_o)
    n141_q <= n140_o;
  initial
    n141_q = 8'b11111111;
  /* vlm5030_gl.vhd:319:7  */
  assign n142_o = n106_o ? 1'b1 : rstdel_block_npor;
  /* vlm5030_gl.vhd:319:7  */
  always @(posedge n103_o)
    n143_q <= n142_o;
  initial
    n143_q = 1'b0;
  /* vlm5030_gl.vhd:335:7  */
  assign n144_o = n132_o ? n135_o : rstdel_block_del;
  /* vlm5030_gl.vhd:335:7  */
  always @(posedge n130_o)
    n145_q <= n144_o;
  initial
    n145_q = 2'b00;
  /* vlm5030_gl.vhd:349:12  */
  always @*
    dq_block_rstq = n207_q; // (isignal)
  initial
    dq_block_rstq = 1'b0;
  /* vlm5030_gl.vhd:350:12  */
  assign dq_block_rstclk = n159_o; // (signal)
  /* vlm5030_gl.vhd:351:12  */
  assign dq_block_ldq = n209_q; // (signal)
  /* vlm5030_gl.vhd:352:12  */
  always @*
    dq_block_maskdq53m = n211_q; // (isignal)
  initial
    dq_block_maskdq53m = 1'b0;
  /* vlm5030_gl.vhd:352:23  */
  always @*
    dq_block_maskdq53s = n213_q; // (isignal)
  initial
    dq_block_maskdq53s = 1'b0;
  assign n150_o = osc[0];
  /* vlm5030_gl.vhd:362:28  */
  assign n154_o = osc[0];
  /* vlm5030_gl.vhd:364:24  */
  assign n155_o = ~dq_block_rstq;
  /* vlm5030_gl.vhd:364:33  */
  assign n156_o = n155_o & rst;
  /* vlm5030_gl.vhd:365:37  */
  assign n157_o = ~rst;
  /* vlm5030_gl.vhd:365:33  */
  assign n158_o = dq_block_rstq & n157_o;
  assign n159_o = {n158_o, n156_o, dq_block_rstq, n154_o};
  assign n166_o = dq_block_rstclk[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n168_o = dq_block_rstclk[3];
  assign n178_o = enpitchlat[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n180_o = enpitchlat[2];
  assign n192_o = enpitchlat[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n194_o = enpitchlat[3];
  assign n202_o = dq_block_ldq[5:3];
  /* vlm5030_gl.vhd:395:7  */
  assign n203_o = maskdq53 ? 3'b000 : n202_o;
  assign n204_o = dq_block_ldq[7:6];
  assign n205_o = dq_block_ldq[2:0];
  /* vlm5030_gl.vhd:357:7  */
  always @(posedge n150_o)
    n207_q <= rst;
  initial
    n207_q = 1'b0;
  /* vlm5030_gl.vhd:369:7  */
  assign n208_o = n168_o ? i_d : dq_block_ldq;
  /* vlm5030_gl.vhd:369:7  */
  always @(posedge n166_o)
    n209_q <= n208_o;
  /* vlm5030_gl.vhd:378:7  */
  assign n210_o = n180_o ? rfdo97zero : dq_block_maskdq53m;
  /* vlm5030_gl.vhd:378:7  */
  always @(posedge n178_o or posedge startrise)
    if (startrise)
      n211_q <= 1'b1;
    else
      n211_q <= n210_o;
  /* vlm5030_gl.vhd:386:7  */
  assign n212_o = n194_o ? dq_block_maskdq53m : dq_block_maskdq53s;
  /* vlm5030_gl.vhd:386:7  */
  always @(posedge n192_o or posedge startrise)
    if (startrise)
      n213_q <= 1'b1;
    else
      n213_q <= n212_o;
  /* vlm5030_gl.vhd:420:12  */
  assign tst_block_ntst1 = n214_o; // (signal)
  /* vlm5030_gl.vhd:420:19  */
  assign tst_block_nstart = n215_o; // (signal)
  /* vlm5030_gl.vhd:420:27  */
  assign tst_block_nvcu = n216_o; // (signal)
  /* vlm5030_gl.vhd:421:12  */
  assign tst_block_ntst1vref = n218_o; // (signal)
  /* vlm5030_gl.vhd:423:15  */
  assign n214_o = ~i_tst1;
  /* vlm5030_gl.vhd:424:15  */
  assign n215_o = ~i_start;
  /* vlm5030_gl.vhd:425:15  */
  assign n216_o = ~i_vcu;
  /* vlm5030_gl.vhd:427:24  */
  assign n217_o = ~(tst_block_nstart | i_tst1);
  /* vlm5030_gl.vhd:429:25  */
  assign n218_o = ~(i_tst1 & i_vref);
  /* vlm5030_gl.vhd:431:31  */
  assign n219_o = tst_block_ntst1 | i_vref;
  /* vlm5030_gl.vhd:431:41  */
  assign n220_o = n219_o | tst_block_nvcu;
  /* vlm5030_gl.vhd:431:50  */
  assign n221_o = n220_o | tst_block_nstart;
  /* vlm5030_gl.vhd:431:20  */
  assign n222_o = ~n221_o;
  /* vlm5030_gl.vhd:432:41  */
  assign n223_o = tst_block_ntst1vref | tst_block_nvcu;
  /* vlm5030_gl.vhd:432:50  */
  assign n224_o = n223_o | i_start;
  /* vlm5030_gl.vhd:432:20  */
  assign n225_o = ~n224_o;
  /* vlm5030_gl.vhd:433:41  */
  assign n226_o = tst_block_ntst1vref | i_vcu;
  /* vlm5030_gl.vhd:433:50  */
  assign n227_o = n226_o | i_start;
  /* vlm5030_gl.vhd:433:20  */
  assign n228_o = ~n227_o;
  /* vlm5030_gl.vhd:433:63  */
  assign n229_o = n228_o | tstenie2dac;
  /* vlm5030_gl.vhd:434:41  */
  assign n230_o = tst_block_ntst1vref | tst_block_nvcu;
  /* vlm5030_gl.vhd:434:50  */
  assign n231_o = n230_o | tst_block_nstart;
  /* vlm5030_gl.vhd:434:20  */
  assign n232_o = ~n231_o;
  /* vlm5030_gl.vhd:435:41  */
  assign n233_o = tst_block_ntst1vref | i_vcu;
  /* vlm5030_gl.vhd:435:50  */
  assign n234_o = n233_o | tst_block_nstart;
  /* vlm5030_gl.vhd:435:20  */
  assign n235_o = ~n234_o;
  /* vlm5030_gl.vhd:436:31  */
  assign n236_o = tst_block_ntst1 | i_vref;
  /* vlm5030_gl.vhd:436:41  */
  assign n237_o = n236_o | i_vcu;
  /* vlm5030_gl.vhd:436:50  */
  assign n238_o = n237_o | tst_block_nstart;
  /* vlm5030_gl.vhd:436:20  */
  assign n239_o = ~n238_o;
  /* vlm5030_gl.vhd:437:31  */
  assign n240_o = tst_block_ntst1 | i_vref;
  /* vlm5030_gl.vhd:437:50  */
  assign n241_o = n240_o | i_start;
  /* vlm5030_gl.vhd:437:20  */
  assign n242_o = ~n241_o;
  /* vlm5030_gl.vhd:448:22  */
  assign n243_o = osc[0];
  assign n251_o = osc[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n253_o = osc[2];
  /* vlm5030_gl.vhd:457:32  */
  assign n256_o = clk2[1];
  /* vlm5030_gl.vhd:457:23  */
  assign n257_o = ~n256_o;
  /* vlm5030_gl.vhd:453:9  */
  assign n258_o = tststopclk2 ? 1'b0 : n257_o;
  /* vlm5030_gl.vhd:462:22  */
  assign n263_o = tststopclk2 ? 1'b0 : n272_o;
  /* vlm5030_gl.vhd:463:22  */
  assign n264_o = osc[2];
  /* clock_functions_pack.vhd:175:17  */
  assign n270_o = clk2[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n271_o = ~n270_o;
  /* vlm5030_gl.vhd:462:45  */
  assign n272_o = n271_o ? n264_o : 1'b0;
  /* vlm5030_gl.vhd:465:22  */
  assign n275_o = tststopclk2 ? 1'b0 : n283_o;
  /* vlm5030_gl.vhd:466:22  */
  assign n276_o = osc[2];
  /* clock_functions_pack.vhd:175:17  */
  assign n282_o = clk2[1];
  /* vlm5030_gl.vhd:465:45  */
  assign n283_o = n282_o ? n276_o : 1'b0;
  /* clock_functions_pack.vhd:75:25  */
  assign n290_o = clk2[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n291_o = clk2[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n292_o = ~n291_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n293_o = clk2[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n294_o = clk2[2];
  assign n295_o = {n294_o, n293_o, n292_o, n290_o};
  /* vlm5030_gl.vhd:479:12  */
  assign clk2div_block_c2qnor = n340_o; // (signal)
  /* vlm5030_gl.vhd:480:12  */
  assign clk2div_block_feedback = n342_o; // (signal)
  assign n303_o = clk2[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n305_o = clk2[2];
  /* vlm5030_gl.vhd:496:29  */
  assign n307_o = clk2divq[9:0];
  /* vlm5030_gl.vhd:496:42  */
  assign n308_o = {n307_o, clk2div_block_feedback};
  /* vlm5030_gl.vhd:500:28  */
  assign n312_o = clk2divq[9:0];
  /* vlm5030_pack.vhd:40:24  */
  assign n318_o = n312_o[9];
  /* vlm5030_pack.vhd:40:20  */
  assign n320_o = 1'b0 | n318_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n322_o = n312_o[8];
  /* vlm5030_pack.vhd:40:20  */
  assign n323_o = n320_o | n322_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n324_o = n312_o[7];
  /* vlm5030_pack.vhd:40:20  */
  assign n325_o = n323_o | n324_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n326_o = n312_o[6];
  /* vlm5030_pack.vhd:40:20  */
  assign n327_o = n325_o | n326_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n328_o = n312_o[5];
  /* vlm5030_pack.vhd:40:20  */
  assign n329_o = n327_o | n328_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n330_o = n312_o[4];
  /* vlm5030_pack.vhd:40:20  */
  assign n331_o = n329_o | n330_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n332_o = n312_o[3];
  /* vlm5030_pack.vhd:40:20  */
  assign n333_o = n331_o | n332_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n334_o = n312_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n335_o = n333_o | n334_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n336_o = n312_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n337_o = n335_o | n336_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n338_o = n312_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n339_o = n337_o | n338_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n340_o = ~n339_o;
  /* vlm5030_gl.vhd:503:21  */
  assign n342_o = rstdel ? 1'b0 : clk2div_block_c2qnor;
  /* vlm5030_gl.vhd:505:64  */
  assign n344_o = clk2divq[0];
  /* vlm5030_gl.vhd:485:30  */
  assign n349_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n350_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n351_o = ~n344_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n352_o = n350_o & n351_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n353_o = n352_o & clk2div_block_feedback;
  /* vlm5030_gl.vhd:488:30  */
  assign n354_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n355_o = n354_o & n344_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n356_o = ~clk2div_block_feedback;
  /* vlm5030_gl.vhd:488:47  */
  assign n357_o = n355_o & n356_o;
  assign n358_o = {n357_o, n353_o, n344_o, n349_o};
  /* vlm5030_gl.vhd:506:64  */
  assign n360_o = clk2divq[1];
  /* vlm5030_gl.vhd:506:88  */
  assign n361_o = clk2divq[0];
  /* vlm5030_gl.vhd:485:30  */
  assign n366_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n367_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n368_o = ~n360_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n369_o = n367_o & n368_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n370_o = n369_o & n361_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n371_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n372_o = n371_o & n360_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n373_o = ~n361_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n374_o = n372_o & n373_o;
  assign n375_o = {n374_o, n370_o, n360_o, n366_o};
  /* vlm5030_gl.vhd:508:64  */
  assign n377_o = clk2divq[3];
  /* vlm5030_gl.vhd:508:88  */
  assign n378_o = clk2divq[2];
  /* vlm5030_gl.vhd:485:30  */
  assign n383_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n384_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n385_o = ~n377_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n386_o = n384_o & n385_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n387_o = n386_o & n378_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n388_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n389_o = n388_o & n377_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n390_o = ~n378_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n391_o = n389_o & n390_o;
  assign n392_o = {n391_o, n387_o, n377_o, n383_o};
  /* vlm5030_gl.vhd:509:64  */
  assign n394_o = clk2divq[4];
  /* vlm5030_gl.vhd:509:88  */
  assign n395_o = clk2divq[3];
  /* vlm5030_gl.vhd:485:30  */
  assign n400_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n401_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n402_o = ~n394_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n403_o = n401_o & n402_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n404_o = n403_o & n395_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n405_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n406_o = n405_o & n394_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n407_o = ~n395_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n408_o = n406_o & n407_o;
  assign n409_o = {n408_o, n404_o, n394_o, n400_o};
  /* vlm5030_gl.vhd:510:64  */
  assign n411_o = clk2divq[5];
  /* vlm5030_gl.vhd:510:88  */
  assign n412_o = clk2divq[4];
  /* vlm5030_gl.vhd:485:30  */
  assign n417_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n418_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n419_o = ~n411_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n420_o = n418_o & n419_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n421_o = n420_o & n412_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n422_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n423_o = n422_o & n411_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n424_o = ~n412_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n425_o = n423_o & n424_o;
  assign n426_o = {n425_o, n421_o, n411_o, n417_o};
  /* vlm5030_gl.vhd:511:64  */
  assign n428_o = clk2divq[6];
  /* vlm5030_gl.vhd:511:88  */
  assign n429_o = clk2divq[5];
  /* vlm5030_gl.vhd:485:30  */
  assign n434_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n435_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n436_o = ~n428_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n437_o = n435_o & n436_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n438_o = n437_o & n429_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n439_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n440_o = n439_o & n428_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n441_o = ~n429_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n442_o = n440_o & n441_o;
  assign n443_o = {n442_o, n438_o, n428_o, n434_o};
  /* vlm5030_gl.vhd:512:64  */
  assign n445_o = clk2divq[7];
  /* vlm5030_gl.vhd:512:88  */
  assign n446_o = clk2divq[6];
  /* vlm5030_gl.vhd:485:30  */
  assign n451_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n452_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n453_o = ~n445_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n454_o = n452_o & n453_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n455_o = n454_o & n446_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n456_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n457_o = n456_o & n445_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n458_o = ~n446_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n459_o = n457_o & n458_o;
  assign n460_o = {n459_o, n455_o, n445_o, n451_o};
  /* vlm5030_gl.vhd:513:64  */
  assign n462_o = clk2divq[8];
  /* vlm5030_gl.vhd:513:88  */
  assign n463_o = clk2divq[7];
  /* vlm5030_gl.vhd:485:30  */
  assign n468_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n469_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n470_o = ~n462_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n471_o = n469_o & n470_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n472_o = n471_o & n463_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n473_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n474_o = n473_o & n462_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n475_o = ~n463_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n476_o = n474_o & n475_o;
  assign n477_o = {n476_o, n472_o, n462_o, n468_o};
  /* vlm5030_gl.vhd:514:64  */
  assign n479_o = clk2divq[9];
  /* vlm5030_gl.vhd:514:88  */
  assign n480_o = clk2divq[8];
  /* vlm5030_gl.vhd:485:30  */
  assign n485_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n486_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n487_o = ~n479_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n488_o = n486_o & n487_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n489_o = n488_o & n480_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n490_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n491_o = n490_o & n479_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n492_o = ~n480_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n493_o = n491_o & n492_o;
  assign n494_o = {n493_o, n489_o, n479_o, n485_o};
  /* vlm5030_gl.vhd:515:64  */
  assign n496_o = clk2divq[10];
  /* vlm5030_gl.vhd:515:88  */
  assign n497_o = clk2divq[9];
  /* vlm5030_gl.vhd:485:30  */
  assign n502_o = clk2[0];
  /* vlm5030_gl.vhd:487:30  */
  assign n503_o = clk2[2];
  /* vlm5030_gl.vhd:487:39  */
  assign n504_o = ~n496_o;
  /* vlm5030_gl.vhd:487:35  */
  assign n505_o = n503_o & n504_o;
  /* vlm5030_gl.vhd:487:47  */
  assign n506_o = n505_o & n497_o;
  /* vlm5030_gl.vhd:488:30  */
  assign n507_o = clk2[2];
  /* vlm5030_gl.vhd:488:35  */
  assign n508_o = n507_o & n496_o;
  /* vlm5030_gl.vhd:488:51  */
  assign n509_o = ~n497_o;
  /* vlm5030_gl.vhd:488:47  */
  assign n510_o = n508_o & n509_o;
  assign n511_o = {n510_o, n506_o, n496_o, n502_o};
  /* vlm5030_gl.vhd:519:5  */
  vlm5030_srlatchclk clk2div_block_c2d5fin_b (
    .i_clk_base(n512_o),
    .i_clk_val(n513_o),
    .i_clk_rise(n514_o),
    .i_clk_fall(n515_o),
    .i_res_base(n516_o),
    .i_res_val(n517_o),
    .i_res_rise(n518_o),
    .i_res_fall(n519_o),
    .i_set_base(n520_o),
    .i_set_val(n521_o),
    .i_set_rise(n522_o),
    .i_set_fall(n523_o),
    .o_q_base(clk2div_block_c2d5fin_b_o_q_base),
    .o_q_val(clk2div_block_c2d5fin_b_o_q_val),
    .o_q_rise(clk2div_block_c2d5fin_b_o_q_rise),
    .o_q_fall(clk2div_block_c2d5fin_b_o_q_fall));
  assign n512_o = osc[0];
  assign n513_o = osc[1];
  assign n514_o = osc[2];
  assign n515_o = osc[3];
  assign n516_o = c2d0[0];
  assign n517_o = c2d0[1];
  assign n518_o = c2d0[2];
  assign n519_o = c2d0[3];
  assign n520_o = c2d5[0];
  assign n521_o = c2d5[1];
  assign n522_o = c2d5[2];
  assign n523_o = c2d5[3];
  assign n524_o = {clk2div_block_c2d5fin_b_o_q_fall, clk2div_block_c2d5fin_b_o_q_rise, clk2div_block_c2d5fin_b_o_q_val, clk2div_block_c2d5fin_b_o_q_base};
  /* vlm5030_gl.vhd:526:5  */
  vlm5030_srlatchclk clk2div_block_c2d7fin_b (
    .i_clk_base(n526_o),
    .i_clk_val(n527_o),
    .i_clk_rise(n528_o),
    .i_clk_fall(n529_o),
    .i_res_base(n530_o),
    .i_res_val(n531_o),
    .i_res_rise(n532_o),
    .i_res_fall(n533_o),
    .i_set_base(n534_o),
    .i_set_val(n535_o),
    .i_set_rise(n536_o),
    .i_set_fall(n537_o),
    .o_q_base(clk2div_block_c2d7fin_b_o_q_base),
    .o_q_val(clk2div_block_c2d7fin_b_o_q_val),
    .o_q_rise(clk2div_block_c2d7fin_b_o_q_rise),
    .o_q_fall(clk2div_block_c2d7fin_b_o_q_fall));
  assign n526_o = osc[0];
  assign n527_o = osc[1];
  assign n528_o = osc[2];
  assign n529_o = osc[3];
  assign n530_o = c2d0[0];
  assign n531_o = c2d0[1];
  assign n532_o = c2d0[2];
  assign n533_o = c2d0[3];
  assign n534_o = c2d7[0];
  assign n535_o = c2d7[1];
  assign n536_o = c2d7[2];
  assign n537_o = c2d7[3];
  assign n538_o = {clk2div_block_c2d7fin_b_o_q_fall, clk2div_block_c2d7fin_b_o_q_rise, clk2div_block_c2d7fin_b_o_q_val, clk2div_block_c2d7fin_b_o_q_base};
  /* clock_functions_pack.vhd:75:25  */
  assign n545_o = c2d7fin[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n546_o = c2d7fin[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n547_o = ~n546_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n548_o = c2d7fin[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n549_o = c2d7fin[2];
  assign n550_o = {n549_o, n548_o, n547_o, n545_o};
  /* vlm5030_gl.vhd:535:5  */
  vlm5030_srlatchclk clk2div_block_c2d9fin_b (
    .i_clk_base(n551_o),
    .i_clk_val(n552_o),
    .i_clk_rise(n553_o),
    .i_clk_fall(n554_o),
    .i_res_base(n555_o),
    .i_res_val(n556_o),
    .i_res_rise(n557_o),
    .i_res_fall(n558_o),
    .i_set_base(n559_o),
    .i_set_val(n560_o),
    .i_set_rise(n561_o),
    .i_set_fall(n562_o),
    .o_q_base(clk2div_block_c2d9fin_b_o_q_base),
    .o_q_val(clk2div_block_c2d9fin_b_o_q_val),
    .o_q_rise(clk2div_block_c2d9fin_b_o_q_rise),
    .o_q_fall(clk2div_block_c2d9fin_b_o_q_fall));
  assign n551_o = osc[0];
  assign n552_o = osc[1];
  assign n553_o = osc[2];
  assign n554_o = osc[3];
  assign n555_o = c2d0[0];
  assign n556_o = c2d0[1];
  assign n557_o = c2d0[2];
  assign n558_o = c2d0[3];
  assign n559_o = c2d9[0];
  assign n560_o = c2d9[1];
  assign n561_o = c2d9[2];
  assign n562_o = c2d9[3];
  assign n563_o = {clk2div_block_c2d9fin_b_o_q_fall, clk2div_block_c2d9fin_b_o_q_rise, clk2div_block_c2d9fin_b_o_q_val, clk2div_block_c2d9fin_b_o_q_base};
  /* clock_functions_pack.vhd:75:25  */
  assign n570_o = c2d9fin[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n571_o = c2d9fin[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n572_o = ~n571_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n573_o = c2d9fin[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n574_o = c2d9fin[2];
  assign n575_o = {n574_o, n573_o, n572_o, n570_o};
  /* clock_functions_pack.vhd:83:26  */
  assign n582_o = c2d5[0];
  /* clock_functions_pack.vhd:84:26  */
  assign n583_o = c2d5[1];
  /* clock_functions_pack.vhd:84:39  */
  assign n584_o = nclk2[1];
  /* clock_functions_pack.vhd:84:30  */
  assign n585_o = n583_o & n584_o;
  /* clock_functions_pack.vhd:85:27  */
  assign n586_o = c2d5[2];
  /* clock_functions_pack.vhd:85:41  */
  assign n587_o = nclk2[1];
  /* clock_functions_pack.vhd:85:32  */
  assign n588_o = n586_o & n587_o;
  /* clock_functions_pack.vhd:85:58  */
  assign n589_o = nclk2[3];
  /* clock_functions_pack.vhd:85:49  */
  assign n590_o = ~n589_o;
  /* clock_functions_pack.vhd:85:45  */
  assign n591_o = n588_o & n590_o;
  /* clock_functions_pack.vhd:86:27  */
  assign n592_o = nclk2[2];
  /* clock_functions_pack.vhd:86:41  */
  assign n593_o = c2d5[1];
  /* clock_functions_pack.vhd:86:32  */
  assign n594_o = n592_o & n593_o;
  /* clock_functions_pack.vhd:86:58  */
  assign n595_o = c2d5[3];
  /* clock_functions_pack.vhd:86:49  */
  assign n596_o = ~n595_o;
  /* clock_functions_pack.vhd:86:45  */
  assign n597_o = n594_o & n596_o;
  /* clock_functions_pack.vhd:85:64  */
  assign n598_o = n591_o | n597_o;
  /* clock_functions_pack.vhd:87:27  */
  assign n599_o = c2d5[3];
  /* clock_functions_pack.vhd:87:41  */
  assign n600_o = nclk2[1];
  /* clock_functions_pack.vhd:87:32  */
  assign n601_o = n599_o & n600_o;
  /* clock_functions_pack.vhd:88:27  */
  assign n602_o = nclk2[3];
  /* clock_functions_pack.vhd:88:41  */
  assign n603_o = c2d5[1];
  /* clock_functions_pack.vhd:88:32  */
  assign n604_o = n602_o & n603_o;
  /* clock_functions_pack.vhd:87:46  */
  assign n605_o = n601_o | n604_o;
  assign n606_o = {n605_o, n598_o, n585_o, n582_o};
  /* clock_functions_pack.vhd:152:26  */
  assign n611_o = c2d0[0];
  /* clock_functions_pack.vhd:153:26  */
  assign n612_o = c2d0[1];
  /* clock_functions_pack.vhd:153:39  */
  assign n613_o = n606_o[1];
  /* clock_functions_pack.vhd:153:30  */
  assign n614_o = ~(n612_o | n613_o);
  /* clock_functions_pack.vhd:154:27  */
  assign n615_o = c2d0[3];
  /* clock_functions_pack.vhd:154:45  */
  assign n616_o = n606_o[1];
  /* clock_functions_pack.vhd:154:36  */
  assign n617_o = ~n616_o;
  /* clock_functions_pack.vhd:154:32  */
  assign n618_o = n615_o & n617_o;
  /* clock_functions_pack.vhd:154:62  */
  assign n619_o = n606_o[2];
  /* clock_functions_pack.vhd:154:53  */
  assign n620_o = ~n619_o;
  /* clock_functions_pack.vhd:154:49  */
  assign n621_o = n618_o & n620_o;
  /* clock_functions_pack.vhd:155:27  */
  assign n622_o = n606_o[3];
  /* clock_functions_pack.vhd:155:45  */
  assign n623_o = c2d0[1];
  /* clock_functions_pack.vhd:155:36  */
  assign n624_o = ~n623_o;
  /* clock_functions_pack.vhd:155:32  */
  assign n625_o = n622_o & n624_o;
  /* clock_functions_pack.vhd:155:62  */
  assign n626_o = c2d0[2];
  /* clock_functions_pack.vhd:155:53  */
  assign n627_o = ~n626_o;
  /* clock_functions_pack.vhd:155:49  */
  assign n628_o = n625_o & n627_o;
  /* clock_functions_pack.vhd:154:68  */
  assign n629_o = n621_o | n628_o;
  /* clock_functions_pack.vhd:156:27  */
  assign n630_o = c2d0[2];
  /* clock_functions_pack.vhd:156:45  */
  assign n631_o = n606_o[1];
  /* clock_functions_pack.vhd:156:36  */
  assign n632_o = ~n631_o;
  /* clock_functions_pack.vhd:156:32  */
  assign n633_o = n630_o & n632_o;
  /* clock_functions_pack.vhd:157:27  */
  assign n634_o = n606_o[2];
  /* clock_functions_pack.vhd:157:45  */
  assign n635_o = c2d0[1];
  /* clock_functions_pack.vhd:157:36  */
  assign n636_o = ~n635_o;
  /* clock_functions_pack.vhd:157:32  */
  assign n637_o = n634_o & n636_o;
  /* clock_functions_pack.vhd:156:50  */
  assign n638_o = n633_o | n637_o;
  assign n639_o = {n638_o, n629_o, n614_o, n611_o};
  /* clock_functions_pack.vhd:75:25  */
  assign n645_o = c2d1[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n646_o = c2d1[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n647_o = ~n646_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n648_o = c2d1[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n649_o = c2d1[2];
  assign n650_o = {n649_o, n648_o, n647_o, n645_o};
  /* clock_functions_pack.vhd:75:25  */
  assign n657_o = c2d3[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n658_o = c2d3[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n659_o = ~n658_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n660_o = c2d3[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n661_o = c2d3[2];
  assign n662_o = {n661_o, n660_o, n659_o, n657_o};
  /* clock_functions_pack.vhd:162:26  */
  assign n667_o = n662_o[0];
  /* clock_functions_pack.vhd:163:26  */
  assign n668_o = n662_o[1];
  /* clock_functions_pack.vhd:163:30  */
  assign n669_o = ~(n668_o | c2d3gate);
  /* clock_functions_pack.vhd:164:26  */
  assign n670_o = n662_o[3];
  /* clock_functions_pack.vhd:164:35  */
  assign n671_o = ~c2d3gate;
  /* clock_functions_pack.vhd:164:31  */
  assign n672_o = n670_o & n671_o;
  /* clock_functions_pack.vhd:165:26  */
  assign n673_o = n662_o[2];
  /* clock_functions_pack.vhd:165:35  */
  assign n674_o = ~c2d3gate;
  /* clock_functions_pack.vhd:165:31  */
  assign n675_o = n673_o & n674_o;
  assign n676_o = {n675_o, n672_o, n669_o, n667_o};
  /* clock_functions_pack.vhd:75:25  */
  assign n682_o = c2d6[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n683_o = c2d6[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n684_o = ~n683_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n685_o = c2d6[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n686_o = c2d6[2];
  assign n687_o = {n686_o, n685_o, n684_o, n682_o};
  /* clock_functions_pack.vhd:75:25  */
  assign n693_o = c2d8[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n694_o = c2d8[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n695_o = ~n694_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n696_o = c2d8[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n697_o = c2d8[2];
  assign n698_o = {n697_o, n696_o, n695_o, n693_o};
  /* clock_functions_pack.vhd:75:25  */
  assign n704_o = c2d10[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n705_o = c2d10[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n706_o = ~n705_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n707_o = c2d10[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n708_o = c2d10[2];
  assign n709_o = {n708_o, n707_o, n706_o, n704_o};
  /* vlm5030_gl.vhd:558:12  */
  assign fsrom_block_fsroma = n1998_q; // (signal)
  assign n717_o = clk2ena[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n719_o = clk2ena[2];
  /* vlm5030_gl.vhd:566:27  */
  assign n721_o = ~(fsromnorlow & nvcufinal);
  /* vlm5030_gl.vhd:566:43  */
  assign n722_o = ~n721_o;
  /* vlm5030_gl.vhd:568:29  */
  assign n723_o = fsrom_block_fsroma[4:0];
  /* vlm5030_gl.vhd:568:51  */
  assign n724_o = fsrom_block_fsroma[0];
  /* vlm5030_gl.vhd:568:65  */
  assign n725_o = fsrom_block_fsroma[5];
  /* vlm5030_gl.vhd:568:55  */
  assign n726_o = n724_o ^ n725_o;
  /* vlm5030_gl.vhd:568:42  */
  assign n727_o = {n723_o, n726_o};
  /* vlm5030_gl.vhd:571:29  */
  assign n728_o = ~rstdel;
  assign n734_o = {1'b0, 1'b0, n728_o, 1'b0};
  assign n735_o = {1'b0, 1'b0};
  assign n736_o = {n734_o, n735_o};
  /* vlm5030_gl.vhd:566:11  */
  assign n737_o = n722_o ? n727_o : n736_o;
  /* vlm5030_gl.vhd:578:38  */
  assign n740_o = fsromdo[9];
  /* vlm5030_gl.vhd:578:54  */
  assign n741_o = xromdo[0];
  /* vlm5030_gl.vhd:578:67  */
  assign n742_o = xromdo[4];
  /* vlm5030_gl.vhd:578:58  */
  assign n743_o = n741_o | n742_o;
  /* vlm5030_gl.vhd:578:43  */
  assign n744_o = n740_o & n743_o;
  /* vlm5030_gl.vhd:579:38  */
  assign n745_o = fsromdo[10];
  /* vlm5030_gl.vhd:579:54  */
  assign n746_o = xromdo[1];
  /* vlm5030_gl.vhd:579:67  */
  assign n747_o = xromdo[4];
  /* vlm5030_gl.vhd:579:58  */
  assign n748_o = n746_o | n747_o;
  /* vlm5030_gl.vhd:579:43  */
  assign n749_o = n745_o & n748_o;
  /* vlm5030_gl.vhd:579:27  */
  assign n750_o = n744_o | n749_o;
  /* vlm5030_gl.vhd:580:38  */
  assign n751_o = fsromdo[11];
  /* vlm5030_gl.vhd:580:54  */
  assign n752_o = xromdo[6];
  /* vlm5030_gl.vhd:580:67  */
  assign n753_o = xromdo[3];
  /* vlm5030_gl.vhd:580:58  */
  assign n754_o = n752_o | n753_o;
  /* vlm5030_gl.vhd:580:80  */
  assign n755_o = xromdo[0];
  /* vlm5030_gl.vhd:580:71  */
  assign n756_o = n754_o | n755_o;
  /* vlm5030_gl.vhd:580:43  */
  assign n757_o = n751_o & n756_o;
  /* vlm5030_gl.vhd:580:27  */
  assign n758_o = n750_o | n757_o;
  /* vlm5030_gl.vhd:581:38  */
  assign n759_o = fsromdo[12];
  /* vlm5030_gl.vhd:581:54  */
  assign n760_o = xromdo[5];
  /* vlm5030_gl.vhd:581:67  */
  assign n761_o = xromdo[2];
  /* vlm5030_gl.vhd:581:58  */
  assign n762_o = n760_o | n761_o;
  /* vlm5030_gl.vhd:581:43  */
  assign n763_o = n759_o & n762_o;
  /* vlm5030_gl.vhd:581:27  */
  assign n764_o = n758_o | n763_o;
  /* vlm5030_gl.vhd:582:38  */
  assign n765_o = fsromdo[13];
  /* vlm5030_gl.vhd:582:54  */
  assign n766_o = xromdo[5];
  /* vlm5030_gl.vhd:582:43  */
  assign n767_o = n765_o & n766_o;
  /* vlm5030_gl.vhd:582:27  */
  assign n768_o = n764_o | n767_o;
  /* vlm5030_gl.vhd:583:38  */
  assign n769_o = fsromdo[8];
  /* vlm5030_gl.vhd:583:54  */
  assign n770_o = xromdo[7];
  /* vlm5030_gl.vhd:583:67  */
  assign n771_o = xromdo[1];
  /* vlm5030_gl.vhd:583:58  */
  assign n772_o = n770_o | n771_o;
  /* vlm5030_gl.vhd:583:43  */
  assign n773_o = n769_o & n772_o;
  /* vlm5030_gl.vhd:583:27  */
  assign n774_o = n768_o | n773_o;
  /* vlm5030_gl.vhd:578:23  */
  assign n775_o = ~n774_o;
  /* vlm5030_gl.vhd:588:14  */
  assign fsrom_block_rom_block_na = n776_o; // (signal)
  /* vlm5030_gl.vhd:589:14  */
  assign fsrom_block_rom_block_ndq = n778_o; // (signal)
  /* vlm5030_gl.vhd:592:14  */
  assign fsrom_block_rom_block_wl = n813_o; // (signal)
  /* vlm5030_gl.vhd:595:14  */
  assign n776_o = ~fsrom_block_fsroma;
  /* vlm5030_gl.vhd:596:20  */
  assign n777_o = dq[5:3];
  /* vlm5030_gl.vhd:596:14  */
  assign n778_o = ~n777_o;
  /* vlm5030_gl.vhd:602:14  */
  assign n779_o = fsrom_block_fsroma[5];
  /* vlm5030_gl.vhd:602:20  */
  assign n780_o = fsrom_block_rom_block_na[5];
  /* vlm5030_gl.vhd:602:17  */
  assign n781_o = {n779_o, n780_o};
  /* vlm5030_gl.vhd:602:28  */
  assign n782_o = fsrom_block_rom_block_na[4];
  /* vlm5030_gl.vhd:602:24  */
  assign n783_o = {n781_o, n782_o};
  /* vlm5030_gl.vhd:602:33  */
  assign n784_o = fsrom_block_fsroma[4];
  /* vlm5030_gl.vhd:602:31  */
  assign n785_o = {n783_o, n784_o};
  /* vlm5030_gl.vhd:602:40  */
  assign n786_o = fsrom_block_fsroma[3];
  /* vlm5030_gl.vhd:602:37  */
  assign n787_o = {n785_o, n786_o};
  /* vlm5030_gl.vhd:602:46  */
  assign n788_o = fsrom_block_rom_block_na[3];
  /* vlm5030_gl.vhd:602:43  */
  assign n789_o = {n787_o, n788_o};
  /* vlm5030_gl.vhd:602:54  */
  assign n790_o = fsrom_block_rom_block_na[2];
  /* vlm5030_gl.vhd:602:50  */
  assign n791_o = {n789_o, n790_o};
  /* vlm5030_gl.vhd:602:59  */
  assign n792_o = fsrom_block_fsroma[2];
  /* vlm5030_gl.vhd:602:57  */
  assign n793_o = {n791_o, n792_o};
  /* vlm5030_gl.vhd:602:66  */
  assign n794_o = fsrom_block_fsroma[1];
  /* vlm5030_gl.vhd:602:63  */
  assign n795_o = {n793_o, n794_o};
  /* vlm5030_gl.vhd:602:72  */
  assign n796_o = fsrom_block_rom_block_na[1];
  /* vlm5030_gl.vhd:602:69  */
  assign n797_o = {n795_o, n796_o};
  /* vlm5030_gl.vhd:602:80  */
  assign n798_o = fsrom_block_rom_block_na[0];
  /* vlm5030_gl.vhd:602:76  */
  assign n799_o = {n797_o, n798_o};
  /* vlm5030_gl.vhd:602:85  */
  assign n800_o = fsrom_block_fsroma[0];
  /* vlm5030_gl.vhd:602:83  */
  assign n801_o = {n799_o, n800_o};
  /* vlm5030_gl.vhd:602:93  */
  assign n802_o = dq[3];
  /* vlm5030_gl.vhd:602:89  */
  assign n803_o = {n801_o, n802_o};
  /* vlm5030_gl.vhd:602:100  */
  assign n804_o = fsrom_block_rom_block_ndq[0];
  /* vlm5030_gl.vhd:602:96  */
  assign n805_o = {n803_o, n804_o};
  /* vlm5030_gl.vhd:602:109  */
  assign n806_o = fsrom_block_rom_block_ndq[1];
  /* vlm5030_gl.vhd:602:104  */
  assign n807_o = {n805_o, n806_o};
  /* vlm5030_gl.vhd:602:115  */
  assign n808_o = dq[4];
  /* vlm5030_gl.vhd:602:112  */
  assign n809_o = {n807_o, n808_o};
  /* vlm5030_gl.vhd:602:123  */
  assign n810_o = dq[5];
  /* vlm5030_gl.vhd:602:119  */
  assign n811_o = {n809_o, n810_o};
  /* vlm5030_gl.vhd:602:130  */
  assign n812_o = fsrom_block_rom_block_ndq[2];
  /* vlm5030_gl.vhd:602:126  */
  assign n813_o = {n811_o, n812_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n820_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n822_o = n820_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n824_o = 1'b0 | n822_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n826_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n828_o = n826_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n829_o = n824_o | n828_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n830_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n832_o = n830_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n833_o = n829_o | n832_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n834_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n836_o = n834_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n837_o = n833_o | n836_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n838_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n840_o = n838_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n841_o = n837_o | n840_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n842_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n844_o = n842_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n845_o = n841_o | n844_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n846_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n848_o = n846_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n849_o = n845_o | n848_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n850_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n852_o = n850_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n853_o = n849_o | n852_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n854_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n856_o = n854_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n857_o = n853_o | n856_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n858_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n860_o = n858_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n861_o = n857_o | n860_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n862_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n864_o = n862_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n865_o = n861_o | n864_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n866_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n868_o = n866_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n869_o = n865_o | n868_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n870_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n872_o = n870_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n873_o = n869_o | n872_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n874_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n876_o = n874_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n877_o = n873_o | n876_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n878_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n880_o = n878_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n881_o = n877_o | n880_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n882_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n884_o = n882_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n885_o = n881_o | n884_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n886_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n888_o = n886_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n889_o = n885_o | n888_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n890_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n892_o = n890_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n893_o = n889_o | n892_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n894_o = ~n893_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n901_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n903_o = n901_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n905_o = 1'b0 | n903_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n907_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n909_o = n907_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n910_o = n905_o | n909_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n911_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n913_o = n911_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n914_o = n910_o | n913_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n915_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n917_o = n915_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n918_o = n914_o | n917_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n919_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n921_o = n919_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n922_o = n918_o | n921_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n923_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n925_o = n923_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n926_o = n922_o | n925_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n927_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n929_o = n927_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n930_o = n926_o | n929_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n931_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n933_o = n931_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n934_o = n930_o | n933_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n935_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n937_o = n935_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n938_o = n934_o | n937_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n939_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n941_o = n939_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n942_o = n938_o | n941_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n943_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n945_o = n943_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n946_o = n942_o | n945_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n947_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n949_o = n947_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n950_o = n946_o | n949_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n951_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n953_o = n951_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n954_o = n950_o | n953_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n955_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n957_o = n955_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n958_o = n954_o | n957_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n959_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n961_o = n959_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n962_o = n958_o | n961_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n963_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n965_o = n963_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n966_o = n962_o | n965_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n967_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n969_o = n967_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n970_o = n966_o | n969_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n971_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n973_o = n971_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n974_o = n970_o | n973_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n975_o = ~n974_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n982_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n984_o = n982_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n986_o = 1'b0 | n984_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n988_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n990_o = n988_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n991_o = n986_o | n990_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n992_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n994_o = n992_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n995_o = n991_o | n994_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n996_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n998_o = n996_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n999_o = n995_o | n998_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1000_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1002_o = n1000_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1003_o = n999_o | n1002_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1004_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1006_o = n1004_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1007_o = n1003_o | n1006_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1008_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1010_o = n1008_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1011_o = n1007_o | n1010_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1012_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1014_o = n1012_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1015_o = n1011_o | n1014_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1016_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1018_o = n1016_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1019_o = n1015_o | n1018_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1020_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1022_o = n1020_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1023_o = n1019_o | n1022_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1024_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1026_o = n1024_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1027_o = n1023_o | n1026_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1028_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1030_o = n1028_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1031_o = n1027_o | n1030_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1032_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1034_o = n1032_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1035_o = n1031_o | n1034_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1036_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1038_o = n1036_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1039_o = n1035_o | n1038_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1040_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1042_o = n1040_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1043_o = n1039_o | n1042_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1044_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1046_o = n1044_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1047_o = n1043_o | n1046_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1048_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1050_o = n1048_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1051_o = n1047_o | n1050_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1052_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1054_o = n1052_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1055_o = n1051_o | n1054_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1056_o = ~n1055_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1063_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1065_o = n1063_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1067_o = 1'b0 | n1065_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1069_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1071_o = n1069_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1072_o = n1067_o | n1071_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1073_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1075_o = n1073_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1076_o = n1072_o | n1075_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1077_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1079_o = n1077_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1080_o = n1076_o | n1079_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1081_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1083_o = n1081_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1084_o = n1080_o | n1083_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1085_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1087_o = n1085_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1088_o = n1084_o | n1087_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1089_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1091_o = n1089_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1092_o = n1088_o | n1091_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1093_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1095_o = n1093_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1096_o = n1092_o | n1095_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1097_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1099_o = n1097_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1100_o = n1096_o | n1099_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1101_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1103_o = n1101_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1104_o = n1100_o | n1103_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1105_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1107_o = n1105_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1108_o = n1104_o | n1107_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1109_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1111_o = n1109_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1112_o = n1108_o | n1111_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1113_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1115_o = n1113_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1116_o = n1112_o | n1115_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1117_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1119_o = n1117_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1120_o = n1116_o | n1119_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1121_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1123_o = n1121_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1124_o = n1120_o | n1123_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1125_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1127_o = n1125_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1128_o = n1124_o | n1127_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1129_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1131_o = n1129_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1132_o = n1128_o | n1131_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1133_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1135_o = n1133_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1136_o = n1132_o | n1135_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1137_o = ~n1136_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1144_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1146_o = n1144_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1148_o = 1'b0 | n1146_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1150_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1152_o = n1150_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1153_o = n1148_o | n1152_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1154_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1156_o = n1154_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1157_o = n1153_o | n1156_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1158_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1160_o = n1158_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1161_o = n1157_o | n1160_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1162_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1164_o = n1162_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1165_o = n1161_o | n1164_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1166_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1168_o = n1166_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1169_o = n1165_o | n1168_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1170_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1172_o = n1170_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1173_o = n1169_o | n1172_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1174_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1176_o = n1174_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1177_o = n1173_o | n1176_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1178_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1180_o = n1178_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1181_o = n1177_o | n1180_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1182_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1184_o = n1182_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1185_o = n1181_o | n1184_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1186_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1188_o = n1186_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1189_o = n1185_o | n1188_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1190_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1192_o = n1190_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1193_o = n1189_o | n1192_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1194_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1196_o = n1194_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1197_o = n1193_o | n1196_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1198_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1200_o = n1198_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1201_o = n1197_o | n1200_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1202_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1204_o = n1202_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1205_o = n1201_o | n1204_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1206_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1208_o = n1206_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1209_o = n1205_o | n1208_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1210_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1212_o = n1210_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1213_o = n1209_o | n1212_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1214_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1216_o = n1214_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1217_o = n1213_o | n1216_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1218_o = ~n1217_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1225_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1227_o = n1225_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1229_o = 1'b0 | n1227_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1231_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1233_o = n1231_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1234_o = n1229_o | n1233_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1235_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1237_o = n1235_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1238_o = n1234_o | n1237_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1239_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1241_o = n1239_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1242_o = n1238_o | n1241_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1243_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1245_o = n1243_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1246_o = n1242_o | n1245_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1247_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1249_o = n1247_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1250_o = n1246_o | n1249_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1251_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1253_o = n1251_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1254_o = n1250_o | n1253_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1255_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1257_o = n1255_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1258_o = n1254_o | n1257_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1259_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1261_o = n1259_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1262_o = n1258_o | n1261_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1263_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1265_o = n1263_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1266_o = n1262_o | n1265_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1267_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1269_o = n1267_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1270_o = n1266_o | n1269_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1271_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1273_o = n1271_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1274_o = n1270_o | n1273_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1275_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1277_o = n1275_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1278_o = n1274_o | n1277_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1279_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1281_o = n1279_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1282_o = n1278_o | n1281_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1283_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1285_o = n1283_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1286_o = n1282_o | n1285_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1287_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1289_o = n1287_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1290_o = n1286_o | n1289_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1291_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1293_o = n1291_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1294_o = n1290_o | n1293_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1295_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1297_o = n1295_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1298_o = n1294_o | n1297_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1299_o = ~n1298_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1306_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1308_o = n1306_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1310_o = 1'b0 | n1308_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1312_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1314_o = n1312_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1315_o = n1310_o | n1314_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1316_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1318_o = n1316_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1319_o = n1315_o | n1318_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1320_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1322_o = n1320_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1323_o = n1319_o | n1322_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1324_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1326_o = n1324_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1327_o = n1323_o | n1326_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1328_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1330_o = n1328_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1331_o = n1327_o | n1330_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1332_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1334_o = n1332_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1335_o = n1331_o | n1334_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1336_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1338_o = n1336_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1339_o = n1335_o | n1338_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1340_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1342_o = n1340_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1343_o = n1339_o | n1342_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1344_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1346_o = n1344_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1347_o = n1343_o | n1346_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1348_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1350_o = n1348_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1351_o = n1347_o | n1350_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1352_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1354_o = n1352_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1355_o = n1351_o | n1354_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1356_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1358_o = n1356_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1359_o = n1355_o | n1358_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1360_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1362_o = n1360_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1363_o = n1359_o | n1362_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1364_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1366_o = n1364_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1367_o = n1363_o | n1366_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1368_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1370_o = n1368_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1371_o = n1367_o | n1370_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1372_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1374_o = n1372_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1375_o = n1371_o | n1374_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1376_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1378_o = n1376_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1379_o = n1375_o | n1378_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1380_o = ~n1379_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1387_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1389_o = n1387_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1391_o = 1'b0 | n1389_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1393_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1395_o = n1393_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1396_o = n1391_o | n1395_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1397_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1399_o = n1397_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1400_o = n1396_o | n1399_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1401_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1403_o = n1401_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1404_o = n1400_o | n1403_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1405_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1407_o = n1405_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1408_o = n1404_o | n1407_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1409_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1411_o = n1409_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1412_o = n1408_o | n1411_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1413_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1415_o = n1413_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1416_o = n1412_o | n1415_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1417_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1419_o = n1417_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1420_o = n1416_o | n1419_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1421_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1423_o = n1421_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1424_o = n1420_o | n1423_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1425_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1427_o = n1425_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1428_o = n1424_o | n1427_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1429_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1431_o = n1429_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1432_o = n1428_o | n1431_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1433_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1435_o = n1433_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1436_o = n1432_o | n1435_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1437_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1439_o = n1437_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1440_o = n1436_o | n1439_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1441_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1443_o = n1441_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1444_o = n1440_o | n1443_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1445_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1447_o = n1445_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1448_o = n1444_o | n1447_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1449_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1451_o = n1449_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1452_o = n1448_o | n1451_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1453_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1455_o = n1453_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1456_o = n1452_o | n1455_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1457_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1459_o = n1457_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1460_o = n1456_o | n1459_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1461_o = ~n1460_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1468_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1470_o = n1468_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1472_o = 1'b0 | n1470_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1474_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1476_o = n1474_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1477_o = n1472_o | n1476_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1478_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1480_o = n1478_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1481_o = n1477_o | n1480_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1482_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1484_o = n1482_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1485_o = n1481_o | n1484_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1486_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1488_o = n1486_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1489_o = n1485_o | n1488_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1490_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1492_o = n1490_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1493_o = n1489_o | n1492_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1494_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1496_o = n1494_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1497_o = n1493_o | n1496_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1498_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1500_o = n1498_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1501_o = n1497_o | n1500_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1502_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1504_o = n1502_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1505_o = n1501_o | n1504_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1506_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1508_o = n1506_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1509_o = n1505_o | n1508_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1510_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1512_o = n1510_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1513_o = n1509_o | n1512_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1514_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1516_o = n1514_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1517_o = n1513_o | n1516_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1518_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1520_o = n1518_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1521_o = n1517_o | n1520_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1522_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1524_o = n1522_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1525_o = n1521_o | n1524_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1526_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1528_o = n1526_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1529_o = n1525_o | n1528_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1530_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1532_o = n1530_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1533_o = n1529_o | n1532_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1534_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1536_o = n1534_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1537_o = n1533_o | n1536_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1538_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1540_o = n1538_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1541_o = n1537_o | n1540_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1542_o = ~n1541_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1549_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1551_o = n1549_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1553_o = 1'b0 | n1551_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1555_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1557_o = n1555_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1558_o = n1553_o | n1557_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1559_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1561_o = n1559_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1562_o = n1558_o | n1561_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1563_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1565_o = n1563_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1566_o = n1562_o | n1565_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1567_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1569_o = n1567_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1570_o = n1566_o | n1569_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1571_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1573_o = n1571_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1574_o = n1570_o | n1573_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1575_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1577_o = n1575_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1578_o = n1574_o | n1577_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1579_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1581_o = n1579_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1582_o = n1578_o | n1581_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1583_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1585_o = n1583_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1586_o = n1582_o | n1585_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1587_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1589_o = n1587_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1590_o = n1586_o | n1589_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1591_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1593_o = n1591_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1594_o = n1590_o | n1593_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1595_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1597_o = n1595_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1598_o = n1594_o | n1597_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1599_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1601_o = n1599_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1602_o = n1598_o | n1601_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1603_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1605_o = n1603_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1606_o = n1602_o | n1605_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1607_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1609_o = n1607_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1610_o = n1606_o | n1609_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1611_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1613_o = n1611_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1614_o = n1610_o | n1613_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1615_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1617_o = n1615_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1618_o = n1614_o | n1617_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1619_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1621_o = n1619_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1622_o = n1618_o | n1621_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1623_o = ~n1622_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1630_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1632_o = n1630_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1634_o = 1'b0 | n1632_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1636_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1638_o = n1636_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1639_o = n1634_o | n1638_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1640_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1642_o = n1640_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1643_o = n1639_o | n1642_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1644_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1646_o = n1644_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1647_o = n1643_o | n1646_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1648_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1650_o = n1648_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1651_o = n1647_o | n1650_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1652_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1654_o = n1652_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1655_o = n1651_o | n1654_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1656_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1658_o = n1656_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1659_o = n1655_o | n1658_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1660_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1662_o = n1660_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1663_o = n1659_o | n1662_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1664_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1666_o = n1664_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1667_o = n1663_o | n1666_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1668_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1670_o = n1668_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1671_o = n1667_o | n1670_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1672_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1674_o = n1672_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1675_o = n1671_o | n1674_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1676_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1678_o = n1676_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1679_o = n1675_o | n1678_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1680_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1682_o = n1680_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1683_o = n1679_o | n1682_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1684_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1686_o = n1684_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1687_o = n1683_o | n1686_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1688_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1690_o = n1688_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1691_o = n1687_o | n1690_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1692_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1694_o = n1692_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1695_o = n1691_o | n1694_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1696_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1698_o = n1696_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1699_o = n1695_o | n1698_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1700_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1702_o = n1700_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1703_o = n1699_o | n1702_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1704_o = ~n1703_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1711_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1713_o = n1711_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1715_o = 1'b0 | n1713_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1717_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1719_o = n1717_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1720_o = n1715_o | n1719_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1721_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1723_o = n1721_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1724_o = n1720_o | n1723_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1725_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1727_o = n1725_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1728_o = n1724_o | n1727_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1729_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1731_o = n1729_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1732_o = n1728_o | n1731_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1733_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1735_o = n1733_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1736_o = n1732_o | n1735_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1737_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1739_o = n1737_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1740_o = n1736_o | n1739_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1741_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1743_o = n1741_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1744_o = n1740_o | n1743_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1745_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1747_o = n1745_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1748_o = n1744_o | n1747_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1749_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1751_o = n1749_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1752_o = n1748_o | n1751_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1753_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1755_o = n1753_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1756_o = n1752_o | n1755_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1757_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1759_o = n1757_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1760_o = n1756_o | n1759_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1761_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1763_o = n1761_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1764_o = n1760_o | n1763_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1765_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1767_o = n1765_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1768_o = n1764_o | n1767_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1769_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1771_o = n1769_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1772_o = n1768_o | n1771_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1773_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1775_o = n1773_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1776_o = n1772_o | n1775_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1777_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1779_o = n1777_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1780_o = n1776_o | n1779_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1781_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1783_o = n1781_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1784_o = n1780_o | n1783_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1785_o = ~n1784_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1792_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1794_o = n1792_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1796_o = 1'b0 | n1794_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1798_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1800_o = n1798_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1801_o = n1796_o | n1800_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1802_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1804_o = n1802_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1805_o = n1801_o | n1804_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1806_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1808_o = n1806_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1809_o = n1805_o | n1808_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1810_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1812_o = n1810_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1813_o = n1809_o | n1812_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1814_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1816_o = n1814_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1817_o = n1813_o | n1816_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1818_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1820_o = n1818_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1821_o = n1817_o | n1820_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1822_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1824_o = n1822_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1825_o = n1821_o | n1824_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1826_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1828_o = n1826_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1829_o = n1825_o | n1828_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1830_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1832_o = n1830_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1833_o = n1829_o | n1832_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1834_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1836_o = n1834_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1837_o = n1833_o | n1836_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1838_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1840_o = n1838_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1841_o = n1837_o | n1840_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1842_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1844_o = n1842_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1845_o = n1841_o | n1844_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1846_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1848_o = n1846_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1849_o = n1845_o | n1848_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1850_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1852_o = n1850_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1853_o = n1849_o | n1852_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1854_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1856_o = n1854_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1857_o = n1853_o | n1856_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1858_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1860_o = n1858_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1861_o = n1857_o | n1860_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1862_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1864_o = n1862_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1865_o = n1861_o | n1864_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1866_o = ~n1865_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1873_o = fsrom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n1875_o = n1873_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1877_o = 1'b0 | n1875_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1879_o = fsrom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n1881_o = n1879_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1882_o = n1877_o | n1881_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1883_o = fsrom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n1885_o = n1883_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1886_o = n1882_o | n1885_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1887_o = fsrom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n1889_o = n1887_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1890_o = n1886_o | n1889_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1891_o = fsrom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n1893_o = n1891_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1894_o = n1890_o | n1893_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1895_o = fsrom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n1897_o = n1895_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1898_o = n1894_o | n1897_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1899_o = fsrom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n1901_o = n1899_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1902_o = n1898_o | n1901_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1903_o = fsrom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n1905_o = n1903_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1906_o = n1902_o | n1905_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1907_o = fsrom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n1909_o = n1907_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1910_o = n1906_o | n1909_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1911_o = fsrom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n1913_o = n1911_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1914_o = n1910_o | n1913_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1915_o = fsrom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n1917_o = n1915_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n1918_o = n1914_o | n1917_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1919_o = fsrom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n1921_o = n1919_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1922_o = n1918_o | n1921_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1923_o = fsrom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n1925_o = n1923_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1926_o = n1922_o | n1925_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1927_o = fsrom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n1929_o = n1927_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1930_o = n1926_o | n1929_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1931_o = fsrom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n1933_o = n1931_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1934_o = n1930_o | n1933_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1935_o = fsrom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n1937_o = n1935_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1938_o = n1934_o | n1937_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1939_o = fsrom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n1941_o = n1939_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1942_o = n1938_o | n1941_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n1943_o = fsrom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n1945_o = n1943_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n1946_o = n1942_o | n1945_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n1947_o = ~n1946_o;
  assign n1948_o = {n1947_o, n1866_o, n1785_o, n1704_o};
  assign n1949_o = {n1623_o, n1542_o, n1461_o, n1380_o};
  assign n1950_o = {n1299_o, n1218_o, n1137_o, n1056_o};
  assign n1951_o = {n975_o, n894_o};
  assign n1952_o = {n1948_o, n1949_o, n1950_o, n1951_o};
  /* vlm5030_gl.vhd:627:35  */
  assign n1954_o = fsromdo[13:8];
  /* vlm5030_pack.vhd:40:24  */
  assign n1960_o = n1954_o[5];
  /* vlm5030_pack.vhd:40:20  */
  assign n1962_o = 1'b0 | n1960_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1964_o = n1954_o[4];
  /* vlm5030_pack.vhd:40:20  */
  assign n1965_o = n1962_o | n1964_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1966_o = n1954_o[3];
  /* vlm5030_pack.vhd:40:20  */
  assign n1967_o = n1965_o | n1966_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1968_o = n1954_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n1969_o = n1967_o | n1968_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1970_o = n1954_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n1971_o = n1969_o | n1970_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1972_o = n1954_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n1973_o = n1971_o | n1972_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n1974_o = ~n1973_o;
  /* vlm5030_gl.vhd:628:35  */
  assign n1976_o = fsromdo[5:0];
  /* vlm5030_pack.vhd:40:24  */
  assign n1982_o = n1976_o[5];
  /* vlm5030_pack.vhd:40:20  */
  assign n1984_o = 1'b0 | n1982_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1986_o = n1976_o[4];
  /* vlm5030_pack.vhd:40:20  */
  assign n1987_o = n1984_o | n1986_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1988_o = n1976_o[3];
  /* vlm5030_pack.vhd:40:20  */
  assign n1989_o = n1987_o | n1988_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1990_o = n1976_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n1991_o = n1989_o | n1990_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1992_o = n1976_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n1993_o = n1991_o | n1992_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n1994_o = n1976_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n1995_o = n1993_o | n1994_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n1996_o = ~n1995_o;
  /* vlm5030_gl.vhd:565:9  */
  assign n1997_o = n719_o ? n737_o : fsrom_block_fsroma;
  /* vlm5030_gl.vhd:565:9  */
  always @(posedge n717_o)
    n1998_q <= n1997_o;
  /* vlm5030_gl.vhd:639:12  */
  assign seqrom_block_gseqroma = n2067_o; // (signal)
  /* vlm5030_gl.vhd:643:14  */
  assign seqrom_block_agen_block_ncen3 = n2023_o; // (signal)
  /* vlm5030_gl.vhd:646:14  */
  always @*
    seqrom_block_agen_block_seqroma = n2070_q; // (isignal)
  initial
    seqrom_block_agen_block_seqroma = 5'b11110;
  /* clock_functions_pack.vhd:170:25  */
  assign n2005_o = c2d10[1];
  /* clock_functions_pack.vhd:170:16  */
  assign n2006_o = ~(tstenctrl2a | n2005_o);
  /* clock_functions_pack.vhd:139:26  */
  assign n2012_o = clk2[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n2013_o = clk2[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n2014_o = n2013_o | ncen1;
  /* clock_functions_pack.vhd:141:26  */
  assign n2015_o = clk2[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n2016_o = ~ncen1;
  /* clock_functions_pack.vhd:141:31  */
  assign n2017_o = n2015_o & n2016_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n2018_o = clk2[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n2019_o = ~ncen1;
  /* clock_functions_pack.vhd:142:31  */
  assign n2020_o = n2018_o & n2019_o;
  assign n2021_o = {n2020_o, n2017_o, n2014_o, n2012_o};
  /* vlm5030_gl.vhd:653:33  */
  assign n2022_o = xromdo[7];
  /* vlm5030_gl.vhd:653:23  */
  assign n2023_o = ~(rstdel | n2022_o);
  /* vlm5030_gl.vhd:654:16  */
  assign n2024_o = ~seqrom_block_agen_block_ncen3;
  assign n2032_o = clk2ctrl[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n2034_o = clk2ctrl[2];
  /* vlm5030_gl.vhd:663:55  */
  assign n2036_o = xromdo[36];
  /* vlm5030_gl.vhd:663:46  */
  assign n2037_o = cen3 | n2036_o;
  /* vlm5030_gl.vhd:663:75  */
  assign n2038_o = seqrom_block_agen_block_seqroma[4];
  /* vlm5030_gl.vhd:663:94  */
  assign n2039_o = seqrom_block_agen_block_seqroma[1];
  /* vlm5030_gl.vhd:663:83  */
  assign n2040_o = ~n2039_o;
  /* vlm5030_gl.vhd:663:79  */
  assign n2041_o = n2038_o ^ n2040_o;
  /* vlm5030_gl.vhd:663:63  */
  assign n2042_o = ~n2041_o;
  /* vlm5030_gl.vhd:663:60  */
  assign n2043_o = n2037_o | n2042_o;
  /* vlm5030_gl.vhd:663:36  */
  assign n2044_o = ~n2043_o;
  /* vlm5030_gl.vhd:663:32  */
  assign n2045_o = ~(rstdel | n2044_o);
  /* vlm5030_gl.vhd:665:19  */
  assign n2046_o = ~cen3;
  /* vlm5030_gl.vhd:666:38  */
  assign n2047_o = seqrom_block_agen_block_seqroma[0];
  /* vlm5030_gl.vhd:666:27  */
  assign n2048_o = ~n2047_o;
  /* vlm5030_gl.vhd:667:34  */
  assign n2049_o = seqrom_block_agen_block_seqroma[1];
  /* vlm5030_gl.vhd:668:34  */
  assign n2050_o = seqrom_block_agen_block_seqroma[2];
  /* vlm5030_gl.vhd:669:34  */
  assign n2051_o = seqrom_block_agen_block_seqroma[3];
  assign n2052_o = {n2051_o, n2050_o, n2049_o, n2048_o};
  assign n2053_o = seqrom_block_agen_block_seqroma[4:1];
  /* vlm5030_gl.vhd:665:11  */
  assign n2054_o = n2046_o ? n2052_o : n2053_o;
  /* vlm5030_gl.vhd:671:20  */
  assign n2055_o = ~seqrom_block_agen_block_ncen3;
  /* vlm5030_gl.vhd:671:11  */
  assign n2057_o = n2055_o ? 4'b1111 : n2054_o;
  /* vlm5030_gl.vhd:675:30  */
  assign n2058_o = xromdo[7];
  assign n2060_o = {n2057_o, n2045_o};
  /* vlm5030_gl.vhd:680:19  */
  assign n2063_o = ~xromdo7nq;
  /* vlm5030_gl.vhd:682:26  */
  assign n2064_o = seqrom_block_agen_block_seqroma[4:1];
  /* vlm5030_gl.vhd:682:52  */
  assign n2065_o = seqrom_block_agen_block_seqroma[0];
  /* vlm5030_gl.vhd:682:41  */
  assign n2066_o = ~n2065_o;
  /* vlm5030_gl.vhd:682:39  */
  assign n2067_o = {n2064_o, n2066_o};
  /* vlm5030_gl.vhd:684:26  */
  assign n2068_o = ~(i_tst1 | xromdo7nq);
  /* vlm5030_gl.vhd:662:9  */
  assign n2069_o = n2034_o ? n2060_o : seqrom_block_agen_block_seqroma;
  /* vlm5030_gl.vhd:662:9  */
  always @(posedge n2032_o)
    n2070_q <= n2069_o;
  initial
    n2070_q = 5'b11110;
  /* vlm5030_gl.vhd:696:15  */
  assign seqrom_block_rom_block_na = n2071_o; // (signal)
  /* vlm5030_gl.vhd:703:14  */
  assign seqrom_block_rom_block_ny = n5019_o; // (signal)
  /* vlm5030_gl.vhd:706:14  */
  assign seqrom_block_rom_block_xwl = n2094_o; // (signal)
  /* vlm5030_gl.vhd:707:14  */
  assign seqrom_block_rom_block_ywl = n5047_o; // (signal)
  /* vlm5030_gl.vhd:710:13  */
  assign n2071_o = ~seqrom_block_gseqroma;
  assign n2072_o = seqrom_block_gseqroma[0];
  assign n2073_o = seqrom_block_rom_block_na[0];
  /* vlm5030_gl.vhd:716:18  */
  assign n2074_o = {n2073_o, n2072_o};
  assign n2075_o = seqrom_block_gseqroma[1];
  /* vlm5030_gl.vhd:716:23  */
  assign n2076_o = {n2074_o, n2075_o};
  assign n2077_o = seqrom_block_rom_block_na[1];
  /* vlm5030_gl.vhd:716:28  */
  assign n2078_o = {n2076_o, n2077_o};
  assign n2079_o = seqrom_block_rom_block_na[2];
  /* vlm5030_gl.vhd:716:34  */
  assign n2080_o = {n2078_o, n2079_o};
  assign n2081_o = seqrom_block_gseqroma[2];
  /* vlm5030_gl.vhd:716:40  */
  assign n2082_o = {n2080_o, n2081_o};
  assign n2083_o = seqrom_block_gseqroma[3];
  /* vlm5030_gl.vhd:716:45  */
  assign n2084_o = {n2082_o, n2083_o};
  assign n2085_o = seqrom_block_rom_block_na[3];
  /* vlm5030_gl.vhd:716:50  */
  assign n2086_o = {n2084_o, n2085_o};
  assign n2087_o = seqrom_block_rom_block_na[4];
  /* vlm5030_gl.vhd:716:56  */
  assign n2088_o = {n2086_o, n2087_o};
  assign n2089_o = seqrom_block_gseqroma[4];
  /* vlm5030_gl.vhd:716:62  */
  assign n2090_o = {n2088_o, n2089_o};
  assign n2091_o = nc2d9fin[1];
  /* vlm5030_gl.vhd:716:67  */
  assign n2092_o = {n2090_o, n2091_o};
  assign n2093_o = c2d9fin[1];
  /* vlm5030_gl.vhd:716:73  */
  assign n2094_o = {n2092_o, n2093_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n2101_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2103_o = n2101_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2105_o = 1'b0 | n2103_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2107_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2109_o = n2107_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2110_o = n2105_o | n2109_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2111_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2113_o = n2111_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2114_o = n2110_o | n2113_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2115_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2117_o = n2115_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2118_o = n2114_o | n2117_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2119_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2121_o = n2119_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2122_o = n2118_o | n2121_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2123_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2125_o = n2123_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2126_o = n2122_o | n2125_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2127_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2129_o = n2127_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2130_o = n2126_o | n2129_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2131_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2133_o = n2131_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2134_o = n2130_o | n2133_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2135_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2137_o = n2135_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2138_o = n2134_o | n2137_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2139_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2141_o = n2139_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2142_o = n2138_o | n2141_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2143_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2145_o = n2143_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2146_o = n2142_o | n2145_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2147_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2149_o = n2147_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2150_o = n2146_o | n2149_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2151_o = ~n2150_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2158_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2160_o = n2158_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2162_o = 1'b0 | n2160_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2164_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2166_o = n2164_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2167_o = n2162_o | n2166_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2168_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2170_o = n2168_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2171_o = n2167_o | n2170_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2172_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2174_o = n2172_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2175_o = n2171_o | n2174_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2176_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2178_o = n2176_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2179_o = n2175_o | n2178_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2180_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2182_o = n2180_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2183_o = n2179_o | n2182_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2184_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2186_o = n2184_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2187_o = n2183_o | n2186_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2188_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2190_o = n2188_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2191_o = n2187_o | n2190_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2192_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2194_o = n2192_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2195_o = n2191_o | n2194_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2196_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2198_o = n2196_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2199_o = n2195_o | n2198_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2200_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2202_o = n2200_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2203_o = n2199_o | n2202_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2204_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2206_o = n2204_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2207_o = n2203_o | n2206_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2208_o = ~n2207_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2215_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2217_o = n2215_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2219_o = 1'b0 | n2217_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2221_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2223_o = n2221_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2224_o = n2219_o | n2223_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2225_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2227_o = n2225_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2228_o = n2224_o | n2227_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2229_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2231_o = n2229_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2232_o = n2228_o | n2231_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2233_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2235_o = n2233_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2236_o = n2232_o | n2235_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2237_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2239_o = n2237_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2240_o = n2236_o | n2239_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2241_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2243_o = n2241_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2244_o = n2240_o | n2243_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2245_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2247_o = n2245_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2248_o = n2244_o | n2247_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2249_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2251_o = n2249_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2252_o = n2248_o | n2251_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2253_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2255_o = n2253_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2256_o = n2252_o | n2255_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2257_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2259_o = n2257_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2260_o = n2256_o | n2259_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2261_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2263_o = n2261_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2264_o = n2260_o | n2263_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2265_o = ~n2264_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2272_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2274_o = n2272_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2276_o = 1'b0 | n2274_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2278_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2280_o = n2278_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2281_o = n2276_o | n2280_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2282_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2284_o = n2282_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2285_o = n2281_o | n2284_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2286_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2288_o = n2286_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2289_o = n2285_o | n2288_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2290_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2292_o = n2290_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2293_o = n2289_o | n2292_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2294_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2296_o = n2294_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2297_o = n2293_o | n2296_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2298_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2300_o = n2298_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2301_o = n2297_o | n2300_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2302_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2304_o = n2302_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2305_o = n2301_o | n2304_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2306_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2308_o = n2306_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2309_o = n2305_o | n2308_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2310_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2312_o = n2310_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2313_o = n2309_o | n2312_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2314_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2316_o = n2314_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2317_o = n2313_o | n2316_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2318_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2320_o = n2318_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2321_o = n2317_o | n2320_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2322_o = ~n2321_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2329_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2331_o = n2329_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2333_o = 1'b0 | n2331_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2335_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2337_o = n2335_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2338_o = n2333_o | n2337_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2339_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2341_o = n2339_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2342_o = n2338_o | n2341_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2343_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2345_o = n2343_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2346_o = n2342_o | n2345_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2347_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2349_o = n2347_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2350_o = n2346_o | n2349_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2351_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2353_o = n2351_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2354_o = n2350_o | n2353_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2355_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2357_o = n2355_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2358_o = n2354_o | n2357_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2359_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2361_o = n2359_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2362_o = n2358_o | n2361_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2363_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2365_o = n2363_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2366_o = n2362_o | n2365_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2367_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2369_o = n2367_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2370_o = n2366_o | n2369_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2371_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2373_o = n2371_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2374_o = n2370_o | n2373_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2375_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2377_o = n2375_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2378_o = n2374_o | n2377_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2379_o = ~n2378_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2386_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2388_o = n2386_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2390_o = 1'b0 | n2388_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2392_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2394_o = n2392_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2395_o = n2390_o | n2394_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2396_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2398_o = n2396_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2399_o = n2395_o | n2398_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2400_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2402_o = n2400_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2403_o = n2399_o | n2402_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2404_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2406_o = n2404_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2407_o = n2403_o | n2406_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2408_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2410_o = n2408_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2411_o = n2407_o | n2410_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2412_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2414_o = n2412_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2415_o = n2411_o | n2414_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2416_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2418_o = n2416_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2419_o = n2415_o | n2418_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2420_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2422_o = n2420_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2423_o = n2419_o | n2422_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2424_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2426_o = n2424_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2427_o = n2423_o | n2426_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2428_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2430_o = n2428_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2431_o = n2427_o | n2430_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2432_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2434_o = n2432_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2435_o = n2431_o | n2434_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2436_o = ~n2435_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2443_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2445_o = n2443_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2447_o = 1'b0 | n2445_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2449_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2451_o = n2449_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2452_o = n2447_o | n2451_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2453_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2455_o = n2453_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2456_o = n2452_o | n2455_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2457_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2459_o = n2457_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2460_o = n2456_o | n2459_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2461_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2463_o = n2461_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2464_o = n2460_o | n2463_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2465_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2467_o = n2465_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2468_o = n2464_o | n2467_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2469_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2471_o = n2469_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2472_o = n2468_o | n2471_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2473_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2475_o = n2473_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2476_o = n2472_o | n2475_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2477_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2479_o = n2477_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2480_o = n2476_o | n2479_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2481_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2483_o = n2481_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2484_o = n2480_o | n2483_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2485_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2487_o = n2485_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2488_o = n2484_o | n2487_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2489_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2491_o = n2489_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2492_o = n2488_o | n2491_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2493_o = ~n2492_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2500_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2502_o = n2500_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2504_o = 1'b0 | n2502_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2506_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2508_o = n2506_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2509_o = n2504_o | n2508_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2510_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2512_o = n2510_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2513_o = n2509_o | n2512_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2514_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2516_o = n2514_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2517_o = n2513_o | n2516_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2518_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2520_o = n2518_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2521_o = n2517_o | n2520_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2522_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2524_o = n2522_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2525_o = n2521_o | n2524_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2526_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2528_o = n2526_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2529_o = n2525_o | n2528_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2530_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2532_o = n2530_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2533_o = n2529_o | n2532_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2534_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2536_o = n2534_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2537_o = n2533_o | n2536_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2538_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2540_o = n2538_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2541_o = n2537_o | n2540_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2542_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2544_o = n2542_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2545_o = n2541_o | n2544_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2546_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2548_o = n2546_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2549_o = n2545_o | n2548_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2550_o = ~n2549_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2557_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2559_o = n2557_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2561_o = 1'b0 | n2559_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2563_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2565_o = n2563_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2566_o = n2561_o | n2565_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2567_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2569_o = n2567_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2570_o = n2566_o | n2569_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2571_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2573_o = n2571_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2574_o = n2570_o | n2573_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2575_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2577_o = n2575_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2578_o = n2574_o | n2577_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2579_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2581_o = n2579_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2582_o = n2578_o | n2581_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2583_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2585_o = n2583_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2586_o = n2582_o | n2585_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2587_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2589_o = n2587_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2590_o = n2586_o | n2589_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2591_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2593_o = n2591_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2594_o = n2590_o | n2593_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2595_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2597_o = n2595_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2598_o = n2594_o | n2597_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2599_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2601_o = n2599_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2602_o = n2598_o | n2601_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2603_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2605_o = n2603_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2606_o = n2602_o | n2605_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2607_o = ~n2606_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2614_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2616_o = n2614_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2618_o = 1'b0 | n2616_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2620_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2622_o = n2620_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2623_o = n2618_o | n2622_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2624_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2626_o = n2624_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2627_o = n2623_o | n2626_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2628_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2630_o = n2628_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2631_o = n2627_o | n2630_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2632_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2634_o = n2632_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2635_o = n2631_o | n2634_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2636_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2638_o = n2636_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2639_o = n2635_o | n2638_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2640_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2642_o = n2640_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2643_o = n2639_o | n2642_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2644_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2646_o = n2644_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2647_o = n2643_o | n2646_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2648_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2650_o = n2648_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2651_o = n2647_o | n2650_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2652_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2654_o = n2652_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2655_o = n2651_o | n2654_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2656_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2658_o = n2656_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2659_o = n2655_o | n2658_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2660_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2662_o = n2660_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2663_o = n2659_o | n2662_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2664_o = ~n2663_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2671_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2673_o = n2671_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2675_o = 1'b0 | n2673_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2677_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2679_o = n2677_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2680_o = n2675_o | n2679_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2681_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2683_o = n2681_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2684_o = n2680_o | n2683_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2685_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2687_o = n2685_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2688_o = n2684_o | n2687_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2689_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2691_o = n2689_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2692_o = n2688_o | n2691_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2693_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2695_o = n2693_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2696_o = n2692_o | n2695_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2697_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2699_o = n2697_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2700_o = n2696_o | n2699_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2701_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2703_o = n2701_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2704_o = n2700_o | n2703_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2705_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2707_o = n2705_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2708_o = n2704_o | n2707_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2709_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2711_o = n2709_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2712_o = n2708_o | n2711_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2713_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2715_o = n2713_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2716_o = n2712_o | n2715_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2717_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2719_o = n2717_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2720_o = n2716_o | n2719_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2721_o = ~n2720_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2728_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2730_o = n2728_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2732_o = 1'b0 | n2730_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2734_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2736_o = n2734_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2737_o = n2732_o | n2736_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2738_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2740_o = n2738_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2741_o = n2737_o | n2740_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2742_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2744_o = n2742_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2745_o = n2741_o | n2744_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2746_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2748_o = n2746_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2749_o = n2745_o | n2748_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2750_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2752_o = n2750_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2753_o = n2749_o | n2752_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2754_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2756_o = n2754_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2757_o = n2753_o | n2756_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2758_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2760_o = n2758_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2761_o = n2757_o | n2760_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2762_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2764_o = n2762_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2765_o = n2761_o | n2764_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2766_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2768_o = n2766_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2769_o = n2765_o | n2768_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2770_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2772_o = n2770_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2773_o = n2769_o | n2772_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2774_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2776_o = n2774_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2777_o = n2773_o | n2776_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2778_o = ~n2777_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2785_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2787_o = n2785_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2789_o = 1'b0 | n2787_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2791_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2793_o = n2791_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2794_o = n2789_o | n2793_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2795_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2797_o = n2795_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2798_o = n2794_o | n2797_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2799_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2801_o = n2799_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2802_o = n2798_o | n2801_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2803_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2805_o = n2803_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2806_o = n2802_o | n2805_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2807_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2809_o = n2807_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2810_o = n2806_o | n2809_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2811_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2813_o = n2811_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2814_o = n2810_o | n2813_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2815_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2817_o = n2815_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2818_o = n2814_o | n2817_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2819_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2821_o = n2819_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2822_o = n2818_o | n2821_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2823_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2825_o = n2823_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2826_o = n2822_o | n2825_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2827_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2829_o = n2827_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2830_o = n2826_o | n2829_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2831_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2833_o = n2831_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2834_o = n2830_o | n2833_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2835_o = ~n2834_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2842_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2844_o = n2842_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2846_o = 1'b0 | n2844_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2848_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2850_o = n2848_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2851_o = n2846_o | n2850_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2852_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2854_o = n2852_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2855_o = n2851_o | n2854_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2856_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2858_o = n2856_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2859_o = n2855_o | n2858_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2860_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2862_o = n2860_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2863_o = n2859_o | n2862_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2864_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2866_o = n2864_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2867_o = n2863_o | n2866_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2868_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2870_o = n2868_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2871_o = n2867_o | n2870_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2872_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2874_o = n2872_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2875_o = n2871_o | n2874_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2876_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2878_o = n2876_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2879_o = n2875_o | n2878_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2880_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2882_o = n2880_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2883_o = n2879_o | n2882_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2884_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2886_o = n2884_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2887_o = n2883_o | n2886_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2888_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2890_o = n2888_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2891_o = n2887_o | n2890_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2892_o = ~n2891_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2899_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2901_o = n2899_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2903_o = 1'b0 | n2901_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2905_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2907_o = n2905_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2908_o = n2903_o | n2907_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2909_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2911_o = n2909_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2912_o = n2908_o | n2911_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2913_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2915_o = n2913_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2916_o = n2912_o | n2915_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2917_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2919_o = n2917_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2920_o = n2916_o | n2919_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2921_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2923_o = n2921_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2924_o = n2920_o | n2923_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2925_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2927_o = n2925_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2928_o = n2924_o | n2927_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2929_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2931_o = n2929_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2932_o = n2928_o | n2931_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2933_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2935_o = n2933_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2936_o = n2932_o | n2935_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2937_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2939_o = n2937_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2940_o = n2936_o | n2939_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2941_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n2943_o = n2941_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2944_o = n2940_o | n2943_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2945_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n2947_o = n2945_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2948_o = n2944_o | n2947_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n2949_o = ~n2948_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2956_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n2958_o = n2956_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2960_o = 1'b0 | n2958_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2962_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n2964_o = n2962_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2965_o = n2960_o | n2964_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2966_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n2968_o = n2966_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2969_o = n2965_o | n2968_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2970_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n2972_o = n2970_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2973_o = n2969_o | n2972_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2974_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n2976_o = n2974_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2977_o = n2973_o | n2976_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2978_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n2980_o = n2978_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2981_o = n2977_o | n2980_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2982_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n2984_o = n2982_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2985_o = n2981_o | n2984_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2986_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n2988_o = n2986_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2989_o = n2985_o | n2988_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2990_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n2992_o = n2990_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n2993_o = n2989_o | n2992_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2994_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n2996_o = n2994_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n2997_o = n2993_o | n2996_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n2998_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3000_o = n2998_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3001_o = n2997_o | n3000_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3002_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3004_o = n3002_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3005_o = n3001_o | n3004_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3006_o = ~n3005_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3013_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3015_o = n3013_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3017_o = 1'b0 | n3015_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3019_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3021_o = n3019_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3022_o = n3017_o | n3021_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3023_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3025_o = n3023_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3026_o = n3022_o | n3025_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3027_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3029_o = n3027_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3030_o = n3026_o | n3029_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3031_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3033_o = n3031_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3034_o = n3030_o | n3033_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3035_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3037_o = n3035_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3038_o = n3034_o | n3037_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3039_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3041_o = n3039_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3042_o = n3038_o | n3041_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3043_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3045_o = n3043_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3046_o = n3042_o | n3045_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3047_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3049_o = n3047_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3050_o = n3046_o | n3049_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3051_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3053_o = n3051_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3054_o = n3050_o | n3053_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3055_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3057_o = n3055_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3058_o = n3054_o | n3057_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3059_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3061_o = n3059_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3062_o = n3058_o | n3061_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3063_o = ~n3062_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3070_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3072_o = n3070_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3074_o = 1'b0 | n3072_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3076_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3078_o = n3076_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3079_o = n3074_o | n3078_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3080_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3082_o = n3080_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3083_o = n3079_o | n3082_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3084_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3086_o = n3084_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3087_o = n3083_o | n3086_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3088_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3090_o = n3088_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3091_o = n3087_o | n3090_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3092_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3094_o = n3092_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3095_o = n3091_o | n3094_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3096_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3098_o = n3096_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3099_o = n3095_o | n3098_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3100_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3102_o = n3100_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3103_o = n3099_o | n3102_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3104_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3106_o = n3104_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3107_o = n3103_o | n3106_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3108_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3110_o = n3108_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3111_o = n3107_o | n3110_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3112_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3114_o = n3112_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3115_o = n3111_o | n3114_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3116_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3118_o = n3116_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3119_o = n3115_o | n3118_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3120_o = ~n3119_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3127_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3129_o = n3127_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3131_o = 1'b0 | n3129_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3133_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3135_o = n3133_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3136_o = n3131_o | n3135_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3137_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3139_o = n3137_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3140_o = n3136_o | n3139_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3141_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3143_o = n3141_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3144_o = n3140_o | n3143_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3145_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3147_o = n3145_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3148_o = n3144_o | n3147_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3149_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3151_o = n3149_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3152_o = n3148_o | n3151_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3153_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3155_o = n3153_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3156_o = n3152_o | n3155_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3157_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3159_o = n3157_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3160_o = n3156_o | n3159_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3161_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3163_o = n3161_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3164_o = n3160_o | n3163_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3165_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3167_o = n3165_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3168_o = n3164_o | n3167_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3169_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3171_o = n3169_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3172_o = n3168_o | n3171_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3173_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3175_o = n3173_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3176_o = n3172_o | n3175_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3177_o = ~n3176_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3184_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3186_o = n3184_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3188_o = 1'b0 | n3186_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3190_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3192_o = n3190_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3193_o = n3188_o | n3192_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3194_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3196_o = n3194_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3197_o = n3193_o | n3196_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3198_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3200_o = n3198_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3201_o = n3197_o | n3200_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3202_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3204_o = n3202_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3205_o = n3201_o | n3204_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3206_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3208_o = n3206_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3209_o = n3205_o | n3208_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3210_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3212_o = n3210_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3213_o = n3209_o | n3212_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3214_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3216_o = n3214_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3217_o = n3213_o | n3216_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3218_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3220_o = n3218_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3221_o = n3217_o | n3220_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3222_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3224_o = n3222_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3225_o = n3221_o | n3224_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3226_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3228_o = n3226_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3229_o = n3225_o | n3228_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3230_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3232_o = n3230_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3233_o = n3229_o | n3232_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3234_o = ~n3233_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3241_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3243_o = n3241_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3245_o = 1'b0 | n3243_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3247_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3249_o = n3247_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3250_o = n3245_o | n3249_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3251_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3253_o = n3251_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3254_o = n3250_o | n3253_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3255_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3257_o = n3255_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3258_o = n3254_o | n3257_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3259_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3261_o = n3259_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3262_o = n3258_o | n3261_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3263_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3265_o = n3263_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3266_o = n3262_o | n3265_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3267_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3269_o = n3267_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3270_o = n3266_o | n3269_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3271_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3273_o = n3271_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3274_o = n3270_o | n3273_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3275_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3277_o = n3275_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3278_o = n3274_o | n3277_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3279_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3281_o = n3279_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3282_o = n3278_o | n3281_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3283_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3285_o = n3283_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3286_o = n3282_o | n3285_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3287_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3289_o = n3287_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3290_o = n3286_o | n3289_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3291_o = ~n3290_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3298_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3300_o = n3298_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3302_o = 1'b0 | n3300_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3304_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3306_o = n3304_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3307_o = n3302_o | n3306_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3308_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3310_o = n3308_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3311_o = n3307_o | n3310_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3312_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3314_o = n3312_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3315_o = n3311_o | n3314_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3316_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3318_o = n3316_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3319_o = n3315_o | n3318_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3320_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3322_o = n3320_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3323_o = n3319_o | n3322_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3324_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3326_o = n3324_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3327_o = n3323_o | n3326_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3328_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3330_o = n3328_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3331_o = n3327_o | n3330_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3332_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3334_o = n3332_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3335_o = n3331_o | n3334_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3336_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3338_o = n3336_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3339_o = n3335_o | n3338_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3340_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3342_o = n3340_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3343_o = n3339_o | n3342_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3344_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3346_o = n3344_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3347_o = n3343_o | n3346_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3348_o = ~n3347_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3355_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3357_o = n3355_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3359_o = 1'b0 | n3357_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3361_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3363_o = n3361_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3364_o = n3359_o | n3363_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3365_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3367_o = n3365_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3368_o = n3364_o | n3367_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3369_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3371_o = n3369_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3372_o = n3368_o | n3371_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3373_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3375_o = n3373_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3376_o = n3372_o | n3375_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3377_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3379_o = n3377_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3380_o = n3376_o | n3379_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3381_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3383_o = n3381_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3384_o = n3380_o | n3383_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3385_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3387_o = n3385_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3388_o = n3384_o | n3387_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3389_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3391_o = n3389_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3392_o = n3388_o | n3391_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3393_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3395_o = n3393_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3396_o = n3392_o | n3395_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3397_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3399_o = n3397_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3400_o = n3396_o | n3399_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3401_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3403_o = n3401_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3404_o = n3400_o | n3403_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3405_o = ~n3404_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3412_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3414_o = n3412_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3416_o = 1'b0 | n3414_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3418_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3420_o = n3418_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3421_o = n3416_o | n3420_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3422_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3424_o = n3422_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3425_o = n3421_o | n3424_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3426_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3428_o = n3426_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3429_o = n3425_o | n3428_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3430_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3432_o = n3430_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3433_o = n3429_o | n3432_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3434_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3436_o = n3434_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3437_o = n3433_o | n3436_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3438_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3440_o = n3438_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3441_o = n3437_o | n3440_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3442_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3444_o = n3442_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3445_o = n3441_o | n3444_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3446_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3448_o = n3446_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3449_o = n3445_o | n3448_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3450_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3452_o = n3450_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3453_o = n3449_o | n3452_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3454_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3456_o = n3454_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3457_o = n3453_o | n3456_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3458_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3460_o = n3458_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3461_o = n3457_o | n3460_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3462_o = ~n3461_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3469_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3471_o = n3469_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3473_o = 1'b0 | n3471_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3475_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3477_o = n3475_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3478_o = n3473_o | n3477_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3479_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3481_o = n3479_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3482_o = n3478_o | n3481_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3483_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3485_o = n3483_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3486_o = n3482_o | n3485_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3487_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3489_o = n3487_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3490_o = n3486_o | n3489_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3491_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3493_o = n3491_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3494_o = n3490_o | n3493_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3495_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3497_o = n3495_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3498_o = n3494_o | n3497_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3499_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3501_o = n3499_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3502_o = n3498_o | n3501_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3503_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3505_o = n3503_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3506_o = n3502_o | n3505_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3507_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3509_o = n3507_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3510_o = n3506_o | n3509_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3511_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3513_o = n3511_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3514_o = n3510_o | n3513_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3515_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3517_o = n3515_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3518_o = n3514_o | n3517_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3519_o = ~n3518_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3526_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3528_o = n3526_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3530_o = 1'b0 | n3528_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3532_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3534_o = n3532_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3535_o = n3530_o | n3534_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3536_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3538_o = n3536_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3539_o = n3535_o | n3538_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3540_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3542_o = n3540_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3543_o = n3539_o | n3542_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3544_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3546_o = n3544_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3547_o = n3543_o | n3546_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3548_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3550_o = n3548_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3551_o = n3547_o | n3550_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3552_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3554_o = n3552_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3555_o = n3551_o | n3554_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3556_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3558_o = n3556_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3559_o = n3555_o | n3558_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3560_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3562_o = n3560_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3563_o = n3559_o | n3562_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3564_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3566_o = n3564_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3567_o = n3563_o | n3566_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3568_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3570_o = n3568_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3571_o = n3567_o | n3570_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3572_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3574_o = n3572_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3575_o = n3571_o | n3574_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3576_o = ~n3575_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3583_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3585_o = n3583_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3587_o = 1'b0 | n3585_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3589_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3591_o = n3589_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3592_o = n3587_o | n3591_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3593_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3595_o = n3593_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3596_o = n3592_o | n3595_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3597_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3599_o = n3597_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3600_o = n3596_o | n3599_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3601_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3603_o = n3601_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3604_o = n3600_o | n3603_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3605_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3607_o = n3605_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3608_o = n3604_o | n3607_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3609_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3611_o = n3609_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3612_o = n3608_o | n3611_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3613_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3615_o = n3613_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3616_o = n3612_o | n3615_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3617_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3619_o = n3617_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3620_o = n3616_o | n3619_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3621_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3623_o = n3621_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3624_o = n3620_o | n3623_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3625_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3627_o = n3625_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3628_o = n3624_o | n3627_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3629_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3631_o = n3629_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3632_o = n3628_o | n3631_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3633_o = ~n3632_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3640_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3642_o = n3640_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3644_o = 1'b0 | n3642_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3646_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3648_o = n3646_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3649_o = n3644_o | n3648_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3650_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3652_o = n3650_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3653_o = n3649_o | n3652_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3654_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3656_o = n3654_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3657_o = n3653_o | n3656_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3658_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3660_o = n3658_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3661_o = n3657_o | n3660_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3662_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3664_o = n3662_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3665_o = n3661_o | n3664_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3666_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3668_o = n3666_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3669_o = n3665_o | n3668_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3670_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3672_o = n3670_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3673_o = n3669_o | n3672_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3674_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3676_o = n3674_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3677_o = n3673_o | n3676_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3678_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3680_o = n3678_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3681_o = n3677_o | n3680_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3682_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3684_o = n3682_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3685_o = n3681_o | n3684_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3686_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3688_o = n3686_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3689_o = n3685_o | n3688_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3690_o = ~n3689_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3697_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3699_o = n3697_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3701_o = 1'b0 | n3699_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3703_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3705_o = n3703_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3706_o = n3701_o | n3705_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3707_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3709_o = n3707_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3710_o = n3706_o | n3709_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3711_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3713_o = n3711_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3714_o = n3710_o | n3713_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3715_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3717_o = n3715_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3718_o = n3714_o | n3717_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3719_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3721_o = n3719_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3722_o = n3718_o | n3721_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3723_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3725_o = n3723_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3726_o = n3722_o | n3725_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3727_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3729_o = n3727_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3730_o = n3726_o | n3729_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3731_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3733_o = n3731_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3734_o = n3730_o | n3733_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3735_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3737_o = n3735_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3738_o = n3734_o | n3737_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3739_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3741_o = n3739_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3742_o = n3738_o | n3741_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3743_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3745_o = n3743_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3746_o = n3742_o | n3745_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3747_o = ~n3746_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3754_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3756_o = n3754_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3758_o = 1'b0 | n3756_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3760_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3762_o = n3760_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3763_o = n3758_o | n3762_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3764_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3766_o = n3764_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3767_o = n3763_o | n3766_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3768_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3770_o = n3768_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3771_o = n3767_o | n3770_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3772_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3774_o = n3772_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3775_o = n3771_o | n3774_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3776_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3778_o = n3776_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3779_o = n3775_o | n3778_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3780_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3782_o = n3780_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3783_o = n3779_o | n3782_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3784_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3786_o = n3784_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3787_o = n3783_o | n3786_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3788_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3790_o = n3788_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3791_o = n3787_o | n3790_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3792_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3794_o = n3792_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3795_o = n3791_o | n3794_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3796_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3798_o = n3796_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3799_o = n3795_o | n3798_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3800_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3802_o = n3800_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3803_o = n3799_o | n3802_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3804_o = ~n3803_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3811_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3813_o = n3811_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3815_o = 1'b0 | n3813_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3817_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3819_o = n3817_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3820_o = n3815_o | n3819_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3821_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3823_o = n3821_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3824_o = n3820_o | n3823_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3825_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3827_o = n3825_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3828_o = n3824_o | n3827_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3829_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3831_o = n3829_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3832_o = n3828_o | n3831_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3833_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3835_o = n3833_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3836_o = n3832_o | n3835_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3837_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3839_o = n3837_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3840_o = n3836_o | n3839_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3841_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3843_o = n3841_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3844_o = n3840_o | n3843_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3845_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3847_o = n3845_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3848_o = n3844_o | n3847_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3849_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3851_o = n3849_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3852_o = n3848_o | n3851_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3853_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3855_o = n3853_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3856_o = n3852_o | n3855_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3857_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3859_o = n3857_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3860_o = n3856_o | n3859_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3861_o = ~n3860_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3868_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3870_o = n3868_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3872_o = 1'b0 | n3870_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3874_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3876_o = n3874_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3877_o = n3872_o | n3876_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3878_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3880_o = n3878_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3881_o = n3877_o | n3880_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3882_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3884_o = n3882_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3885_o = n3881_o | n3884_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3886_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3888_o = n3886_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3889_o = n3885_o | n3888_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3890_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3892_o = n3890_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3893_o = n3889_o | n3892_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3894_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3896_o = n3894_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3897_o = n3893_o | n3896_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3898_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3900_o = n3898_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3901_o = n3897_o | n3900_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3902_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3904_o = n3902_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3905_o = n3901_o | n3904_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3906_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3908_o = n3906_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3909_o = n3905_o | n3908_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3910_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3912_o = n3910_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3913_o = n3909_o | n3912_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3914_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3916_o = n3914_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3917_o = n3913_o | n3916_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3918_o = ~n3917_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3925_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3927_o = n3925_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3929_o = 1'b0 | n3927_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3931_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3933_o = n3931_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3934_o = n3929_o | n3933_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3935_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3937_o = n3935_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3938_o = n3934_o | n3937_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3939_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3941_o = n3939_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3942_o = n3938_o | n3941_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3943_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n3945_o = n3943_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3946_o = n3942_o | n3945_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3947_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n3949_o = n3947_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3950_o = n3946_o | n3949_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3951_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n3953_o = n3951_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3954_o = n3950_o | n3953_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3955_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n3957_o = n3955_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3958_o = n3954_o | n3957_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3959_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n3961_o = n3959_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3962_o = n3958_o | n3961_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3963_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n3965_o = n3963_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3966_o = n3962_o | n3965_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3967_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n3969_o = n3967_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3970_o = n3966_o | n3969_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3971_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n3973_o = n3971_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3974_o = n3970_o | n3973_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n3975_o = ~n3974_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3982_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n3984_o = n3982_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3986_o = 1'b0 | n3984_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3988_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n3990_o = n3988_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3991_o = n3986_o | n3990_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3992_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n3994_o = n3992_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n3995_o = n3991_o | n3994_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n3996_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n3998_o = n3996_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n3999_o = n3995_o | n3998_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4000_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4002_o = n4000_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4003_o = n3999_o | n4002_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4004_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4006_o = n4004_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4007_o = n4003_o | n4006_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4008_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4010_o = n4008_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4011_o = n4007_o | n4010_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4012_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4014_o = n4012_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4015_o = n4011_o | n4014_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4016_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n4018_o = n4016_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4019_o = n4015_o | n4018_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4020_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n4022_o = n4020_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4023_o = n4019_o | n4022_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4024_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n4026_o = n4024_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4027_o = n4023_o | n4026_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4028_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n4030_o = n4028_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4031_o = n4027_o | n4030_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n4032_o = ~n4031_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4039_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n4041_o = n4039_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4043_o = 1'b0 | n4041_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4045_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n4047_o = n4045_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4048_o = n4043_o | n4047_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4049_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n4051_o = n4049_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4052_o = n4048_o | n4051_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4053_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n4055_o = n4053_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4056_o = n4052_o | n4055_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4057_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4059_o = n4057_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4060_o = n4056_o | n4059_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4061_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4063_o = n4061_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4064_o = n4060_o | n4063_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4065_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4067_o = n4065_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4068_o = n4064_o | n4067_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4069_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4071_o = n4069_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4072_o = n4068_o | n4071_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4073_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n4075_o = n4073_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4076_o = n4072_o | n4075_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4077_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n4079_o = n4077_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4080_o = n4076_o | n4079_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4081_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n4083_o = n4081_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4084_o = n4080_o | n4083_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4085_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n4087_o = n4085_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4088_o = n4084_o | n4087_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n4089_o = ~n4088_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4096_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n4098_o = n4096_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4100_o = 1'b0 | n4098_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4102_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n4104_o = n4102_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4105_o = n4100_o | n4104_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4106_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n4108_o = n4106_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4109_o = n4105_o | n4108_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4110_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n4112_o = n4110_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4113_o = n4109_o | n4112_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4114_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4116_o = n4114_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4117_o = n4113_o | n4116_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4118_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4120_o = n4118_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4121_o = n4117_o | n4120_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4122_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4124_o = n4122_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4125_o = n4121_o | n4124_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4126_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4128_o = n4126_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4129_o = n4125_o | n4128_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4130_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n4132_o = n4130_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4133_o = n4129_o | n4132_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4134_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n4136_o = n4134_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4137_o = n4133_o | n4136_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4138_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n4140_o = n4138_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4141_o = n4137_o | n4140_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4142_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n4144_o = n4142_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4145_o = n4141_o | n4144_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n4146_o = ~n4145_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4153_o = seqrom_block_rom_block_xwl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n4155_o = n4153_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4157_o = 1'b0 | n4155_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4159_o = seqrom_block_rom_block_xwl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n4161_o = n4159_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4162_o = n4157_o | n4161_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4163_o = seqrom_block_rom_block_xwl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n4165_o = n4163_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4166_o = n4162_o | n4165_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4167_o = seqrom_block_rom_block_xwl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n4169_o = n4167_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4170_o = n4166_o | n4169_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4171_o = seqrom_block_rom_block_xwl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4173_o = n4171_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4174_o = n4170_o | n4173_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4175_o = seqrom_block_rom_block_xwl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4177_o = n4175_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4178_o = n4174_o | n4177_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4179_o = seqrom_block_rom_block_xwl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4181_o = n4179_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4182_o = n4178_o | n4181_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4183_o = seqrom_block_rom_block_xwl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4185_o = n4183_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4186_o = n4182_o | n4185_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4187_o = seqrom_block_rom_block_xwl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n4189_o = n4187_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4190_o = n4186_o | n4189_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4191_o = seqrom_block_rom_block_xwl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n4193_o = n4191_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4194_o = n4190_o | n4193_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4195_o = seqrom_block_rom_block_xwl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n4197_o = n4195_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4198_o = n4194_o | n4197_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4199_o = seqrom_block_rom_block_xwl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n4201_o = n4199_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4202_o = n4198_o | n4201_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n4203_o = ~n4202_o;
  assign n4204_o = {n4203_o, n4146_o, n4089_o, n4032_o};
  assign n4205_o = {n3975_o, n3918_o, n3861_o, n3804_o};
  assign n4206_o = {n3747_o, n3690_o, n3633_o, n3576_o};
  assign n4207_o = {n3519_o, n3462_o, n3405_o, n3348_o};
  assign n4208_o = {n3291_o, n3234_o, n3177_o, n3120_o};
  assign n4209_o = {n3063_o, n3006_o, n2949_o, n2892_o};
  assign n4210_o = {n2835_o, n2778_o, n2721_o, n2664_o};
  assign n4211_o = {n2607_o, n2550_o, n2493_o, n2436_o};
  assign n4212_o = {n2379_o, n2322_o, n2265_o, n2208_o};
  assign n4213_o = {n4204_o, n4205_o, n4206_o, n4207_o};
  assign n4214_o = {n4208_o, n4209_o, n4210_o, n4211_o};
  assign n4215_o = {n4212_o, n2151_o};
  assign n4216_o = {n4213_o, n4214_o, n4215_o};
  /* vlm5030_gl.vhd:772:27  */
  assign n4217_o = xromdo[0];
  /* vlm5030_gl.vhd:772:27  */
  assign n4218_o = xromdo[1];
  /* vlm5030_gl.vhd:772:27  */
  assign n4219_o = xromdo[2];
  /* vlm5030_gl.vhd:772:27  */
  assign n4220_o = xromdo[3];
  /* vlm5030_gl.vhd:772:27  */
  assign n4221_o = xromdo[4];
  /* vlm5030_gl.vhd:772:27  */
  assign n4222_o = xromdo[5];
  /* vlm5030_gl.vhd:772:27  */
  assign n4223_o = xromdo[6];
  /* vlm5030_gl.vhd:772:27  */
  assign n4224_o = xromdo[7];
  /* vlm5030_gl.vhd:772:27  */
  assign n4225_o = xromdo[8];
  /* vlm5030_gl.vhd:772:27  */
  assign n4226_o = xromdo[9];
  /* vlm5030_gl.vhd:772:27  */
  assign n4227_o = xromdo[10];
  /* vlm5030_gl.vhd:772:27  */
  assign n4228_o = xromdo[11];
  /* vlm5030_gl.vhd:772:27  */
  assign n4229_o = xromdo[12];
  /* vlm5030_gl.vhd:772:27  */
  assign n4230_o = xromdo[13];
  /* vlm5030_gl.vhd:772:27  */
  assign n4231_o = xromdo[14];
  /* vlm5030_gl.vhd:772:27  */
  assign n4232_o = xromdo[15];
  /* vlm5030_gl.vhd:772:27  */
  assign n4233_o = xromdo[16];
  /* vlm5030_gl.vhd:772:27  */
  assign n4234_o = xromdo[17];
  /* vlm5030_gl.vhd:772:27  */
  assign n4235_o = xromdo[18];
  /* vlm5030_gl.vhd:772:27  */
  assign n4236_o = xromdo[19];
  /* vlm5030_gl.vhd:772:27  */
  assign n4237_o = xromdo[20];
  /* vlm5030_gl.vhd:772:27  */
  assign n4238_o = xromdo[21];
  /* vlm5030_gl.vhd:772:27  */
  assign n4239_o = xromdo[22];
  /* vlm5030_gl.vhd:772:27  */
  assign n4240_o = xromdo[23];
  /* vlm5030_gl.vhd:772:27  */
  assign n4241_o = xromdo[24];
  /* vlm5030_gl.vhd:772:27  */
  assign n4242_o = xromdo[25];
  /* vlm5030_gl.vhd:772:27  */
  assign n4243_o = xromdo[26];
  /* vlm5030_gl.vhd:772:27  */
  assign n4244_o = xromdo[27];
  /* vlm5030_gl.vhd:772:27  */
  assign n4245_o = xromdo[28];
  /* vlm5030_gl.vhd:772:27  */
  assign n4246_o = xromdo[29];
  /* vlm5030_gl.vhd:772:27  */
  assign n4247_o = xromdo[30];
  /* vlm5030_gl.vhd:772:27  */
  assign n4248_o = xromdo[31];
  /* vlm5030_gl.vhd:772:27  */
  assign n4249_o = xromdo[32];
  /* vlm5030_gl.vhd:772:27  */
  assign n4250_o = xromdo[33];
  /* vlm5030_gl.vhd:772:27  */
  assign n4251_o = xromdo[34];
  /* vlm5030_gl.vhd:772:27  */
  assign n4252_o = xromdo[35];
  /* vlm5030_pack.vhd:50:26  */
  assign n4259_o = seqrom_block_rom_block_ywl[35];
  /* vlm5030_pack.vhd:50:32  */
  assign n4261_o = n4259_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4263_o = 1'b0 | n4261_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4265_o = seqrom_block_rom_block_ywl[34];
  /* vlm5030_pack.vhd:50:32  */
  assign n4267_o = n4265_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4268_o = n4263_o | n4267_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4269_o = seqrom_block_rom_block_ywl[33];
  /* vlm5030_pack.vhd:50:32  */
  assign n4271_o = n4269_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4272_o = n4268_o | n4271_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4273_o = seqrom_block_rom_block_ywl[32];
  /* vlm5030_pack.vhd:50:32  */
  assign n4275_o = n4273_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4276_o = n4272_o | n4275_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4277_o = seqrom_block_rom_block_ywl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n4279_o = n4277_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4280_o = n4276_o | n4279_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4281_o = seqrom_block_rom_block_ywl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n4283_o = n4281_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4284_o = n4280_o | n4283_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4285_o = seqrom_block_rom_block_ywl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n4287_o = n4285_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4288_o = n4284_o | n4287_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4289_o = seqrom_block_rom_block_ywl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n4291_o = n4289_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4292_o = n4288_o | n4291_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4293_o = seqrom_block_rom_block_ywl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n4295_o = n4293_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4296_o = n4292_o | n4295_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4297_o = seqrom_block_rom_block_ywl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n4299_o = n4297_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4300_o = n4296_o | n4299_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4301_o = seqrom_block_rom_block_ywl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n4303_o = n4301_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4304_o = n4300_o | n4303_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4305_o = seqrom_block_rom_block_ywl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n4307_o = n4305_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4308_o = n4304_o | n4307_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4309_o = seqrom_block_rom_block_ywl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n4311_o = n4309_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4312_o = n4308_o | n4311_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4313_o = seqrom_block_rom_block_ywl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n4315_o = n4313_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4316_o = n4312_o | n4315_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4317_o = seqrom_block_rom_block_ywl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n4319_o = n4317_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4320_o = n4316_o | n4319_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4321_o = seqrom_block_rom_block_ywl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n4323_o = n4321_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4324_o = n4320_o | n4323_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4325_o = seqrom_block_rom_block_ywl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n4327_o = n4325_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4328_o = n4324_o | n4327_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4329_o = seqrom_block_rom_block_ywl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n4331_o = n4329_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4332_o = n4328_o | n4331_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4333_o = seqrom_block_rom_block_ywl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n4335_o = n4333_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4336_o = n4332_o | n4335_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4337_o = seqrom_block_rom_block_ywl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n4339_o = n4337_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4340_o = n4336_o | n4339_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4341_o = seqrom_block_rom_block_ywl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n4343_o = n4341_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4344_o = n4340_o | n4343_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4345_o = seqrom_block_rom_block_ywl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n4347_o = n4345_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4348_o = n4344_o | n4347_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4349_o = seqrom_block_rom_block_ywl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n4351_o = n4349_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4352_o = n4348_o | n4351_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4353_o = seqrom_block_rom_block_ywl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n4355_o = n4353_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4356_o = n4352_o | n4355_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4357_o = seqrom_block_rom_block_ywl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n4359_o = n4357_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4360_o = n4356_o | n4359_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4361_o = seqrom_block_rom_block_ywl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n4363_o = n4361_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4364_o = n4360_o | n4363_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4365_o = seqrom_block_rom_block_ywl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n4367_o = n4365_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4368_o = n4364_o | n4367_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4369_o = seqrom_block_rom_block_ywl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n4371_o = n4369_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4372_o = n4368_o | n4371_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4373_o = seqrom_block_rom_block_ywl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4375_o = n4373_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4376_o = n4372_o | n4375_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4377_o = seqrom_block_rom_block_ywl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4379_o = n4377_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4380_o = n4376_o | n4379_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4381_o = seqrom_block_rom_block_ywl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4383_o = n4381_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4384_o = n4380_o | n4383_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4385_o = seqrom_block_rom_block_ywl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4387_o = n4385_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4388_o = n4384_o | n4387_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4389_o = seqrom_block_rom_block_ywl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n4391_o = n4389_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4392_o = n4388_o | n4391_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4393_o = seqrom_block_rom_block_ywl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n4395_o = n4393_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4396_o = n4392_o | n4395_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4397_o = seqrom_block_rom_block_ywl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n4399_o = n4397_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4400_o = n4396_o | n4399_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4401_o = seqrom_block_rom_block_ywl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n4403_o = n4401_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4404_o = n4400_o | n4403_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n4405_o = ~n4404_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4412_o = seqrom_block_rom_block_ywl[35];
  /* vlm5030_pack.vhd:50:32  */
  assign n4414_o = n4412_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4416_o = 1'b0 | n4414_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4418_o = seqrom_block_rom_block_ywl[34];
  /* vlm5030_pack.vhd:50:32  */
  assign n4420_o = n4418_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4421_o = n4416_o | n4420_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4422_o = seqrom_block_rom_block_ywl[33];
  /* vlm5030_pack.vhd:50:32  */
  assign n4424_o = n4422_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4425_o = n4421_o | n4424_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4426_o = seqrom_block_rom_block_ywl[32];
  /* vlm5030_pack.vhd:50:32  */
  assign n4428_o = n4426_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4429_o = n4425_o | n4428_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4430_o = seqrom_block_rom_block_ywl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n4432_o = n4430_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4433_o = n4429_o | n4432_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4434_o = seqrom_block_rom_block_ywl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n4436_o = n4434_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4437_o = n4433_o | n4436_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4438_o = seqrom_block_rom_block_ywl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n4440_o = n4438_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4441_o = n4437_o | n4440_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4442_o = seqrom_block_rom_block_ywl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n4444_o = n4442_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4445_o = n4441_o | n4444_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4446_o = seqrom_block_rom_block_ywl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n4448_o = n4446_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4449_o = n4445_o | n4448_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4450_o = seqrom_block_rom_block_ywl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n4452_o = n4450_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4453_o = n4449_o | n4452_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4454_o = seqrom_block_rom_block_ywl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n4456_o = n4454_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4457_o = n4453_o | n4456_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4458_o = seqrom_block_rom_block_ywl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n4460_o = n4458_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4461_o = n4457_o | n4460_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4462_o = seqrom_block_rom_block_ywl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n4464_o = n4462_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4465_o = n4461_o | n4464_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4466_o = seqrom_block_rom_block_ywl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n4468_o = n4466_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4469_o = n4465_o | n4468_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4470_o = seqrom_block_rom_block_ywl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n4472_o = n4470_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4473_o = n4469_o | n4472_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4474_o = seqrom_block_rom_block_ywl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n4476_o = n4474_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4477_o = n4473_o | n4476_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4478_o = seqrom_block_rom_block_ywl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n4480_o = n4478_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4481_o = n4477_o | n4480_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4482_o = seqrom_block_rom_block_ywl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n4484_o = n4482_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4485_o = n4481_o | n4484_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4486_o = seqrom_block_rom_block_ywl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n4488_o = n4486_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4489_o = n4485_o | n4488_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4490_o = seqrom_block_rom_block_ywl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n4492_o = n4490_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4493_o = n4489_o | n4492_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4494_o = seqrom_block_rom_block_ywl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n4496_o = n4494_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4497_o = n4493_o | n4496_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4498_o = seqrom_block_rom_block_ywl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n4500_o = n4498_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4501_o = n4497_o | n4500_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4502_o = seqrom_block_rom_block_ywl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n4504_o = n4502_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4505_o = n4501_o | n4504_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4506_o = seqrom_block_rom_block_ywl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n4508_o = n4506_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4509_o = n4505_o | n4508_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4510_o = seqrom_block_rom_block_ywl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n4512_o = n4510_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4513_o = n4509_o | n4512_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4514_o = seqrom_block_rom_block_ywl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n4516_o = n4514_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4517_o = n4513_o | n4516_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4518_o = seqrom_block_rom_block_ywl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n4520_o = n4518_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4521_o = n4517_o | n4520_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4522_o = seqrom_block_rom_block_ywl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n4524_o = n4522_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4525_o = n4521_o | n4524_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4526_o = seqrom_block_rom_block_ywl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4528_o = n4526_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4529_o = n4525_o | n4528_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4530_o = seqrom_block_rom_block_ywl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4532_o = n4530_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4533_o = n4529_o | n4532_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4534_o = seqrom_block_rom_block_ywl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4536_o = n4534_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4537_o = n4533_o | n4536_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4538_o = seqrom_block_rom_block_ywl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4540_o = n4538_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4541_o = n4537_o | n4540_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4542_o = seqrom_block_rom_block_ywl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n4544_o = n4542_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4545_o = n4541_o | n4544_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4546_o = seqrom_block_rom_block_ywl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n4548_o = n4546_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4549_o = n4545_o | n4548_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4550_o = seqrom_block_rom_block_ywl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n4552_o = n4550_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4553_o = n4549_o | n4552_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4554_o = seqrom_block_rom_block_ywl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n4556_o = n4554_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4557_o = n4553_o | n4556_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n4558_o = ~n4557_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4565_o = seqrom_block_rom_block_ywl[35];
  /* vlm5030_pack.vhd:50:32  */
  assign n4567_o = n4565_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4569_o = 1'b0 | n4567_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4571_o = seqrom_block_rom_block_ywl[34];
  /* vlm5030_pack.vhd:50:32  */
  assign n4573_o = n4571_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4574_o = n4569_o | n4573_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4575_o = seqrom_block_rom_block_ywl[33];
  /* vlm5030_pack.vhd:50:32  */
  assign n4577_o = n4575_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4578_o = n4574_o | n4577_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4579_o = seqrom_block_rom_block_ywl[32];
  /* vlm5030_pack.vhd:50:32  */
  assign n4581_o = n4579_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4582_o = n4578_o | n4581_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4583_o = seqrom_block_rom_block_ywl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n4585_o = n4583_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4586_o = n4582_o | n4585_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4587_o = seqrom_block_rom_block_ywl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n4589_o = n4587_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4590_o = n4586_o | n4589_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4591_o = seqrom_block_rom_block_ywl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n4593_o = n4591_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4594_o = n4590_o | n4593_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4595_o = seqrom_block_rom_block_ywl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n4597_o = n4595_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4598_o = n4594_o | n4597_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4599_o = seqrom_block_rom_block_ywl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n4601_o = n4599_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4602_o = n4598_o | n4601_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4603_o = seqrom_block_rom_block_ywl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n4605_o = n4603_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4606_o = n4602_o | n4605_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4607_o = seqrom_block_rom_block_ywl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n4609_o = n4607_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4610_o = n4606_o | n4609_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4611_o = seqrom_block_rom_block_ywl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n4613_o = n4611_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4614_o = n4610_o | n4613_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4615_o = seqrom_block_rom_block_ywl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n4617_o = n4615_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4618_o = n4614_o | n4617_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4619_o = seqrom_block_rom_block_ywl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n4621_o = n4619_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4622_o = n4618_o | n4621_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4623_o = seqrom_block_rom_block_ywl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n4625_o = n4623_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4626_o = n4622_o | n4625_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4627_o = seqrom_block_rom_block_ywl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n4629_o = n4627_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4630_o = n4626_o | n4629_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4631_o = seqrom_block_rom_block_ywl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n4633_o = n4631_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4634_o = n4630_o | n4633_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4635_o = seqrom_block_rom_block_ywl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n4637_o = n4635_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4638_o = n4634_o | n4637_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4639_o = seqrom_block_rom_block_ywl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n4641_o = n4639_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4642_o = n4638_o | n4641_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4643_o = seqrom_block_rom_block_ywl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n4645_o = n4643_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4646_o = n4642_o | n4645_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4647_o = seqrom_block_rom_block_ywl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n4649_o = n4647_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4650_o = n4646_o | n4649_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4651_o = seqrom_block_rom_block_ywl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n4653_o = n4651_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4654_o = n4650_o | n4653_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4655_o = seqrom_block_rom_block_ywl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n4657_o = n4655_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4658_o = n4654_o | n4657_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4659_o = seqrom_block_rom_block_ywl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n4661_o = n4659_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4662_o = n4658_o | n4661_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4663_o = seqrom_block_rom_block_ywl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n4665_o = n4663_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4666_o = n4662_o | n4665_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4667_o = seqrom_block_rom_block_ywl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n4669_o = n4667_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4670_o = n4666_o | n4669_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4671_o = seqrom_block_rom_block_ywl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n4673_o = n4671_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4674_o = n4670_o | n4673_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4675_o = seqrom_block_rom_block_ywl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n4677_o = n4675_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4678_o = n4674_o | n4677_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4679_o = seqrom_block_rom_block_ywl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4681_o = n4679_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4682_o = n4678_o | n4681_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4683_o = seqrom_block_rom_block_ywl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4685_o = n4683_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4686_o = n4682_o | n4685_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4687_o = seqrom_block_rom_block_ywl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4689_o = n4687_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4690_o = n4686_o | n4689_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4691_o = seqrom_block_rom_block_ywl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4693_o = n4691_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4694_o = n4690_o | n4693_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4695_o = seqrom_block_rom_block_ywl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n4697_o = n4695_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4698_o = n4694_o | n4697_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4699_o = seqrom_block_rom_block_ywl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n4701_o = n4699_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4702_o = n4698_o | n4701_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4703_o = seqrom_block_rom_block_ywl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n4705_o = n4703_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4706_o = n4702_o | n4705_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4707_o = seqrom_block_rom_block_ywl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n4709_o = n4707_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4710_o = n4706_o | n4709_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n4711_o = ~n4710_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4718_o = seqrom_block_rom_block_ywl[35];
  /* vlm5030_pack.vhd:50:32  */
  assign n4720_o = n4718_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4722_o = 1'b0 | n4720_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4724_o = seqrom_block_rom_block_ywl[34];
  /* vlm5030_pack.vhd:50:32  */
  assign n4726_o = n4724_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4727_o = n4722_o | n4726_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4728_o = seqrom_block_rom_block_ywl[33];
  /* vlm5030_pack.vhd:50:32  */
  assign n4730_o = n4728_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4731_o = n4727_o | n4730_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4732_o = seqrom_block_rom_block_ywl[32];
  /* vlm5030_pack.vhd:50:32  */
  assign n4734_o = n4732_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4735_o = n4731_o | n4734_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4736_o = seqrom_block_rom_block_ywl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n4738_o = n4736_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4739_o = n4735_o | n4738_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4740_o = seqrom_block_rom_block_ywl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n4742_o = n4740_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4743_o = n4739_o | n4742_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4744_o = seqrom_block_rom_block_ywl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n4746_o = n4744_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4747_o = n4743_o | n4746_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4748_o = seqrom_block_rom_block_ywl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n4750_o = n4748_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4751_o = n4747_o | n4750_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4752_o = seqrom_block_rom_block_ywl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n4754_o = n4752_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4755_o = n4751_o | n4754_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4756_o = seqrom_block_rom_block_ywl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n4758_o = n4756_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4759_o = n4755_o | n4758_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4760_o = seqrom_block_rom_block_ywl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n4762_o = n4760_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4763_o = n4759_o | n4762_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4764_o = seqrom_block_rom_block_ywl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n4766_o = n4764_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4767_o = n4763_o | n4766_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4768_o = seqrom_block_rom_block_ywl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n4770_o = n4768_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4771_o = n4767_o | n4770_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4772_o = seqrom_block_rom_block_ywl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n4774_o = n4772_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4775_o = n4771_o | n4774_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4776_o = seqrom_block_rom_block_ywl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n4778_o = n4776_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4779_o = n4775_o | n4778_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4780_o = seqrom_block_rom_block_ywl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n4782_o = n4780_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4783_o = n4779_o | n4782_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4784_o = seqrom_block_rom_block_ywl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n4786_o = n4784_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4787_o = n4783_o | n4786_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4788_o = seqrom_block_rom_block_ywl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n4790_o = n4788_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4791_o = n4787_o | n4790_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4792_o = seqrom_block_rom_block_ywl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n4794_o = n4792_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4795_o = n4791_o | n4794_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4796_o = seqrom_block_rom_block_ywl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n4798_o = n4796_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4799_o = n4795_o | n4798_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4800_o = seqrom_block_rom_block_ywl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n4802_o = n4800_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4803_o = n4799_o | n4802_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4804_o = seqrom_block_rom_block_ywl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n4806_o = n4804_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4807_o = n4803_o | n4806_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4808_o = seqrom_block_rom_block_ywl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n4810_o = n4808_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4811_o = n4807_o | n4810_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4812_o = seqrom_block_rom_block_ywl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n4814_o = n4812_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4815_o = n4811_o | n4814_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4816_o = seqrom_block_rom_block_ywl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n4818_o = n4816_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4819_o = n4815_o | n4818_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4820_o = seqrom_block_rom_block_ywl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n4822_o = n4820_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4823_o = n4819_o | n4822_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4824_o = seqrom_block_rom_block_ywl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n4826_o = n4824_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4827_o = n4823_o | n4826_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4828_o = seqrom_block_rom_block_ywl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n4830_o = n4828_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4831_o = n4827_o | n4830_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4832_o = seqrom_block_rom_block_ywl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4834_o = n4832_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4835_o = n4831_o | n4834_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4836_o = seqrom_block_rom_block_ywl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4838_o = n4836_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4839_o = n4835_o | n4838_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4840_o = seqrom_block_rom_block_ywl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4842_o = n4840_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4843_o = n4839_o | n4842_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4844_o = seqrom_block_rom_block_ywl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4846_o = n4844_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4847_o = n4843_o | n4846_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4848_o = seqrom_block_rom_block_ywl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n4850_o = n4848_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4851_o = n4847_o | n4850_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4852_o = seqrom_block_rom_block_ywl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n4854_o = n4852_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4855_o = n4851_o | n4854_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4856_o = seqrom_block_rom_block_ywl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n4858_o = n4856_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4859_o = n4855_o | n4858_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4860_o = seqrom_block_rom_block_ywl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n4862_o = n4860_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4863_o = n4859_o | n4862_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n4864_o = ~n4863_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4871_o = seqrom_block_rom_block_ywl[35];
  /* vlm5030_pack.vhd:50:32  */
  assign n4873_o = n4871_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4875_o = 1'b0 | n4873_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4877_o = seqrom_block_rom_block_ywl[34];
  /* vlm5030_pack.vhd:50:32  */
  assign n4879_o = n4877_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4880_o = n4875_o | n4879_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4881_o = seqrom_block_rom_block_ywl[33];
  /* vlm5030_pack.vhd:50:32  */
  assign n4883_o = n4881_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4884_o = n4880_o | n4883_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4885_o = seqrom_block_rom_block_ywl[32];
  /* vlm5030_pack.vhd:50:32  */
  assign n4887_o = n4885_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4888_o = n4884_o | n4887_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4889_o = seqrom_block_rom_block_ywl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n4891_o = n4889_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4892_o = n4888_o | n4891_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4893_o = seqrom_block_rom_block_ywl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n4895_o = n4893_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4896_o = n4892_o | n4895_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4897_o = seqrom_block_rom_block_ywl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n4899_o = n4897_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4900_o = n4896_o | n4899_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4901_o = seqrom_block_rom_block_ywl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n4903_o = n4901_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4904_o = n4900_o | n4903_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4905_o = seqrom_block_rom_block_ywl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n4907_o = n4905_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4908_o = n4904_o | n4907_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4909_o = seqrom_block_rom_block_ywl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n4911_o = n4909_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4912_o = n4908_o | n4911_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4913_o = seqrom_block_rom_block_ywl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n4915_o = n4913_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4916_o = n4912_o | n4915_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4917_o = seqrom_block_rom_block_ywl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n4919_o = n4917_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4920_o = n4916_o | n4919_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4921_o = seqrom_block_rom_block_ywl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n4923_o = n4921_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4924_o = n4920_o | n4923_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4925_o = seqrom_block_rom_block_ywl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n4927_o = n4925_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4928_o = n4924_o | n4927_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4929_o = seqrom_block_rom_block_ywl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n4931_o = n4929_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4932_o = n4928_o | n4931_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4933_o = seqrom_block_rom_block_ywl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n4935_o = n4933_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4936_o = n4932_o | n4935_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4937_o = seqrom_block_rom_block_ywl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n4939_o = n4937_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4940_o = n4936_o | n4939_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4941_o = seqrom_block_rom_block_ywl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n4943_o = n4941_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4944_o = n4940_o | n4943_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4945_o = seqrom_block_rom_block_ywl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n4947_o = n4945_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4948_o = n4944_o | n4947_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4949_o = seqrom_block_rom_block_ywl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n4951_o = n4949_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4952_o = n4948_o | n4951_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4953_o = seqrom_block_rom_block_ywl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n4955_o = n4953_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4956_o = n4952_o | n4955_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4957_o = seqrom_block_rom_block_ywl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n4959_o = n4957_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4960_o = n4956_o | n4959_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4961_o = seqrom_block_rom_block_ywl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n4963_o = n4961_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4964_o = n4960_o | n4963_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4965_o = seqrom_block_rom_block_ywl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n4967_o = n4965_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4968_o = n4964_o | n4967_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4969_o = seqrom_block_rom_block_ywl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n4971_o = n4969_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n4972_o = n4968_o | n4971_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4973_o = seqrom_block_rom_block_ywl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n4975_o = n4973_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4976_o = n4972_o | n4975_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4977_o = seqrom_block_rom_block_ywl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n4979_o = n4977_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4980_o = n4976_o | n4979_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4981_o = seqrom_block_rom_block_ywl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n4983_o = n4981_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4984_o = n4980_o | n4983_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4985_o = seqrom_block_rom_block_ywl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n4987_o = n4985_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4988_o = n4984_o | n4987_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4989_o = seqrom_block_rom_block_ywl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n4991_o = n4989_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4992_o = n4988_o | n4991_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4993_o = seqrom_block_rom_block_ywl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n4995_o = n4993_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n4996_o = n4992_o | n4995_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n4997_o = seqrom_block_rom_block_ywl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n4999_o = n4997_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5000_o = n4996_o | n4999_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5001_o = seqrom_block_rom_block_ywl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n5003_o = n5001_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5004_o = n5000_o | n5003_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5005_o = seqrom_block_rom_block_ywl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n5007_o = n5005_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5008_o = n5004_o | n5007_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5009_o = seqrom_block_rom_block_ywl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n5011_o = n5009_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5012_o = n5008_o | n5011_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5013_o = seqrom_block_rom_block_ywl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n5015_o = n5013_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5016_o = n5012_o | n5015_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n5017_o = ~n5016_o;
  assign n5018_o = {n4405_o, n4558_o, n4711_o, n4864_o};
  assign n5019_o = {n5018_o, n5017_o};
  /* vlm5030_gl.vhd:789:30  */
  assign n5021_o = xromdo[7:0];
  /* vlm5030_pack.vhd:40:24  */
  assign n5027_o = n5021_o[7];
  /* vlm5030_pack.vhd:40:20  */
  assign n5029_o = 1'b0 | n5027_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5031_o = n5021_o[6];
  /* vlm5030_pack.vhd:40:20  */
  assign n5032_o = n5029_o | n5031_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5033_o = n5021_o[5];
  /* vlm5030_pack.vhd:40:20  */
  assign n5034_o = n5032_o | n5033_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5035_o = n5021_o[4];
  /* vlm5030_pack.vhd:40:20  */
  assign n5036_o = n5034_o | n5035_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5037_o = n5021_o[3];
  /* vlm5030_pack.vhd:40:20  */
  assign n5038_o = n5036_o | n5037_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5039_o = n5021_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n5040_o = n5038_o | n5039_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5041_o = n5021_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n5042_o = n5040_o | n5041_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5043_o = n5021_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n5044_o = n5042_o | n5043_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n5045_o = ~n5044_o;
  /* vlm5030_gl.vhd:791:17  */
  assign n5046_o = ~seqrom_block_rom_block_ny;
  assign n5047_o = {n4217_o, n4218_o, n4219_o, n4220_o, n4221_o, n4222_o, n4223_o, n4224_o, n4225_o, n4226_o, n4227_o, n4228_o, n4229_o, n4230_o, n4231_o, n4232_o, n4233_o, n4234_o, n4235_o, n4236_o, n4237_o, n4238_o, n4239_o, n4240_o, n4241_o, n4242_o, n4243_o, n4244_o, n4245_o, n4246_o, n4247_o, n4248_o, n4249_o, n4250_o, n4251_o, n4252_o};
  /* vlm5030_gl.vhd:805:12  */
  always @*
    cntdown_block_cntq = n5077_q; // (isignal)
  initial
    cntdown_block_cntq = 5'b00000;
  assign n5056_o = clkcntdn[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5058_o = clkcntdn[2];
  /* vlm5030_gl.vhd:810:23  */
  assign n5060_o = ~ncntdnload;
  /* vlm5030_gl.vhd:811:46  */
  assign n5061_o = dinalq[7:4];
  /* vlm5030_gl.vhd:815:21  */
  assign n5063_o = ~ncntdn;
  /* vlm5030_gl.vhd:816:26  */
  assign n5065_o = cntdown_block_cntq - 5'b00001;
  /* vlm5030_gl.vhd:815:11  */
  assign n5066_o = n5063_o ? n5065_o : cntdown_block_cntq;
  assign n5067_o = {n5061_o, 1'b1};
  /* vlm5030_gl.vhd:810:9  */
  assign n5068_o = n5060_o ? n5067_o : n5066_o;
  /* vlm5030_gl.vhd:823:29  */
  assign n5073_o = cntdown_block_cntq == 5'b00000;
  /* vlm5030_gl.vhd:823:19  */
  assign n5074_o = n5073_o ? 1'b1 : 1'b0;
  /* vlm5030_gl.vhd:809:7  */
  assign n5076_o = n5058_o ? n5068_o : cntdown_block_cntq;
  /* vlm5030_gl.vhd:809:7  */
  always @(posedge n5056_o)
    n5077_q <= n5076_o;
  initial
    n5077_q = 5'b00000;
  /* vlm5030_gl.vhd:833:12  */
  always @*
    din_block_dinlat = n5169_q; // (isignal)
  initial
    din_block_dinlat = 8'b00000000;
  /* vlm5030_gl.vhd:834:12  */
  assign din_block_ndincom = n5113_o; // (signal)
  /* vlm5030_gl.vhd:836:12  */
  assign din_block_latchhq = n5171_q; // (signal)
  /* vlm5030_gl.vhd:836:21  */
  assign din_block_latchh = n5172_o; // (signal)
  assign n5081_o = osc[0];
  /* vlm5030_gl.vhd:842:19  */
  assign n5083_o = ~clkdin;
  /* vlm5030_gl.vhd:848:38  */
  assign n5088_o = xromdo[7:0];
  /* vlm5030_gl.vhd:848:28  */
  assign n5089_o = din_block_dinlat & n5088_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5095_o = n5089_o[7];
  /* vlm5030_pack.vhd:40:20  */
  assign n5097_o = 1'b0 | n5095_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5099_o = n5089_o[6];
  /* vlm5030_pack.vhd:40:20  */
  assign n5100_o = n5097_o | n5099_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5101_o = n5089_o[5];
  /* vlm5030_pack.vhd:40:20  */
  assign n5102_o = n5100_o | n5101_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5103_o = n5089_o[4];
  /* vlm5030_pack.vhd:40:20  */
  assign n5104_o = n5102_o | n5103_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5105_o = n5089_o[3];
  /* vlm5030_pack.vhd:40:20  */
  assign n5106_o = n5104_o | n5105_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5107_o = n5089_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n5108_o = n5106_o | n5107_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5109_o = n5089_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n5110_o = n5108_o | n5109_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5111_o = n5089_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n5112_o = n5110_o | n5111_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n5113_o = ~n5112_o;
  assign n5121_o = c2d3gated[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5123_o = c2d3gated[2];
  /* vlm5030_gl.vhd:855:19  */
  assign n5125_o = ~din_block_ndincom;
  /* vlm5030_gl.vhd:855:39  */
  assign n5126_o = dinalq[7:1];
  /* vlm5030_gl.vhd:855:31  */
  assign n5127_o = {n5125_o, n5126_o};
  assign n5134_o = osc[0];
  /* vlm5030_gl.vhd:868:24  */
  assign n5139_o = dinalq[0];
  /* vlm5030_gl.vhd:868:28  */
  assign n5140_o = eavcu ? n5139_o : n5141_o;
  /* vlm5030_gl.vhd:869:25  */
  assign n5141_o = din_block_latchhq[0];
  /* vlm5030_gl.vhd:870:44  */
  assign n5143_o = eavcu ? 7'b0000000 : n5144_o;
  /* vlm5030_gl.vhd:871:35  */
  assign n5144_o = din_block_latchhq[7:1];
  assign n5152_o = clk2ena[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5154_o = clk2ena[2];
  /* vlm5030_gl.vhd:876:20  */
  assign n5156_o = ~neaload;
  /* vlm5030_gl.vhd:878:51  */
  assign n5157_o = dinalq[0];
  /* vlm5030_gl.vhd:878:41  */
  assign n5158_o = ~n5157_o;
  /* vlm5030_gl.vhd:878:36  */
  assign n5159_o = ~(eavcu | n5158_o);
  /* vlm5030_gl.vhd:879:36  */
  assign n5160_o = dinalq[7:1];
  /* vlm5030_gl.vhd:884:49  */
  assign n5162_o = aq + 16'b0000000000000001;
  /* vlm5030_gl.vhd:882:11  */
  assign n5163_o = eainc ? n5162_o : aq;
  assign n5164_o = {din_block_latchh, n5160_o, n5159_o};
  /* vlm5030_gl.vhd:876:9  */
  assign n5165_o = n5156_o ? n5164_o : n5163_o;
  /* vlm5030_gl.vhd:841:7  */
  assign n5168_o = n5083_o ? i_d : din_block_dinlat;
  /* vlm5030_gl.vhd:841:7  */
  always @(posedge n5081_o)
    n5169_q <= n5168_o;
  initial
    n5169_q = 8'b00000000;
  /* vlm5030_gl.vhd:861:7  */
  assign n5170_o = ealatchh ? dinalq : din_block_latchhq;
  /* vlm5030_gl.vhd:861:7  */
  always @(posedge n5134_o)
    n5171_q <= n5170_o;
  /* vlm5030_gl.vhd:861:7  */
  assign n5172_o = {n5143_o, n5140_o};
  /* vlm5030_gl.vhd:898:12  */
  always @*
    random_block_lfsr = n5224_q; // (isignal)
  initial
    random_block_lfsr = 10'b0000000000;
  /* vlm5030_gl.vhd:899:12  */
  assign random_block_all0 = n5201_o; // (signal)
  /* vlm5030_gl.vhd:900:12  */
  assign random_block_feedback = n5205_o; // (signal)
  /* vlm5030_gl.vhd:903:22  */
  assign n5175_o = random_block_lfsr[8:0];
  /* vlm5030_pack.vhd:40:24  */
  assign n5181_o = n5175_o[8];
  /* vlm5030_pack.vhd:40:20  */
  assign n5183_o = 1'b0 | n5181_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5185_o = n5175_o[7];
  /* vlm5030_pack.vhd:40:20  */
  assign n5186_o = n5183_o | n5185_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5187_o = n5175_o[6];
  /* vlm5030_pack.vhd:40:20  */
  assign n5188_o = n5186_o | n5187_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5189_o = n5175_o[5];
  /* vlm5030_pack.vhd:40:20  */
  assign n5190_o = n5188_o | n5189_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5191_o = n5175_o[4];
  /* vlm5030_pack.vhd:40:20  */
  assign n5192_o = n5190_o | n5191_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5193_o = n5175_o[3];
  /* vlm5030_pack.vhd:40:20  */
  assign n5194_o = n5192_o | n5193_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5195_o = n5175_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n5196_o = n5194_o | n5195_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5197_o = n5175_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n5198_o = n5196_o | n5197_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n5199_o = n5175_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n5200_o = n5198_o | n5199_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n5201_o = ~n5200_o;
  /* vlm5030_gl.vhd:905:22  */
  assign n5202_o = random_block_lfsr[9];
  /* vlm5030_gl.vhd:905:34  */
  assign n5203_o = random_block_lfsr[2];
  /* vlm5030_gl.vhd:905:26  */
  assign n5204_o = n5202_o ^ n5203_o;
  /* vlm5030_gl.vhd:905:39  */
  assign n5205_o = ~(n5204_o | random_block_all0);
  assign n5213_o = clk2ena[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5215_o = clk2ena[2];
  /* vlm5030_gl.vhd:910:21  */
  assign n5217_o = random_block_lfsr[8:0];
  /* vlm5030_gl.vhd:910:44  */
  assign n5218_o = ~(rstdel | random_block_feedback);
  /* vlm5030_gl.vhd:910:34  */
  assign n5219_o = {n5217_o, n5218_o};
  /* vlm5030_gl.vhd:914:19  */
  assign n5222_o = random_block_lfsr[9];
  /* vlm5030_gl.vhd:909:7  */
  assign n5223_o = n5215_o ? n5219_o : random_block_lfsr;
  /* vlm5030_gl.vhd:909:7  */
  always @(posedge n5213_o)
    n5224_q <= n5223_o;
  initial
    n5224_q = 10'b0000000000;
  /* vlm5030_gl.vhd:925:12  */
  assign start_block_nvcu = n5233_o; // (signal)
  /* vlm5030_gl.vhd:927:12  */
  assign start_block_startq = n5722_q; // (signal)
  /* vlm5030_gl.vhd:931:12  */
  assign start_block_startriseq = n5724_q; // (signal)
  /* vlm5030_gl.vhd:932:12  */
  assign start_block_startriseqvcu = n5261_o; // (signal)
  /* vlm5030_gl.vhd:934:12  */
  assign start_block_ffsset = n5262_o; // (signal)
  /* vlm5030_gl.vhd:935:12  */
  assign start_block_ffsloop = n5319_o; // (signal)
  /* vlm5030_gl.vhd:936:12  */
  always @*
    start_block_ffs1q = n5726_q; // (isignal)
  initial
    start_block_ffs1q = 1'b1;
  /* vlm5030_gl.vhd:936:19  */
  always @*
    start_block_ffs2q = n5730_q; // (isignal)
  initial
    start_block_ffs2q = 1'b1;
  /* vlm5030_gl.vhd:937:12  */
  always @*
    start_block_ffs3q = n5732_q; // (isignal)
  initial
    start_block_ffs3q = 1'b1;
  /* vlm5030_gl.vhd:937:19  */
  always @*
    start_block_ffs4q = n5734_q; // (isignal)
  initial
    start_block_ffs4q = 1'b1;
  /* vlm5030_gl.vhd:938:12  */
  assign start_block_ffs1nq = n5310_o; // (signal)
  /* vlm5030_gl.vhd:938:20  */
  assign start_block_ffs2nq = n5311_o; // (signal)
  /* vlm5030_gl.vhd:939:12  */
  assign start_block_ffs3nq = n5312_o; // (signal)
  /* vlm5030_gl.vhd:939:20  */
  assign start_block_ffs4nq = n5313_o; // (signal)
  /* vlm5030_gl.vhd:940:12  */
  always @*
    start_block_ffs5q = n5736_q; // (isignal)
  initial
    start_block_ffs5q = 1'b0;
  /* vlm5030_gl.vhd:941:12  */
  assign start_block_ffs5nq = n5314_o; // (signal)
  /* vlm5030_gl.vhd:942:12  */
  assign start_block_vcumode = n5234_o; // (signal)
  /* vlm5030_gl.vhd:945:12  */
  assign start_block_vcufinal = n5235_o; // (signal)
  /* vlm5030_gl.vhd:946:12  */
  assign start_block_vcufinal1q = n5738_q; // (signal)
  /* vlm5030_gl.vhd:947:12  */
  assign start_block_vcufinal2q = n5740_q; // (signal)
  /* vlm5030_gl.vhd:948:12  */
  assign start_block_nvcufinal12 = n5344_o; // (signal)
  /* vlm5030_gl.vhd:950:12  */
  assign start_block_xromdo7nqdel = start_block_xromdo7nqdel_b_o_out; // (signal)
  /* vlm5030_gl.vhd:952:12  */
  always @*
    start_block_msff1q = n5742_q; // (isignal)
  initial
    start_block_msff1q = 1'b0;
  /* vlm5030_gl.vhd:952:20  */
  always @*
    start_block_msff2q = n5744_q; // (isignal)
  initial
    start_block_msff2q = 1'b0;
  /* vlm5030_gl.vhd:953:12  */
  always @*
    start_block_pmsff3q = n5746_q; // (isignal)
  initial
    start_block_pmsff3q = 1'b0;
  /* vlm5030_gl.vhd:954:12  */
  assign start_block_msff1nq = n5388_o; // (signal)
  /* vlm5030_gl.vhd:954:21  */
  assign start_block_msff2nq = n5408_o; // (signal)
  /* vlm5030_gl.vhd:955:12  */
  assign start_block_pmsff3nq = n5426_o; // (signal)
  /* vlm5030_gl.vhd:956:12  */
  assign start_block_msffset = n5369_o; // (signal)
  /* vlm5030_gl.vhd:958:12  */
  assign start_block_n001x = n5432_o; // (signal)
  /* vlm5030_gl.vhd:958:19  */
  assign start_block_n002x = n5436_o; // (signal)
  /* vlm5030_gl.vhd:958:26  */
  assign start_block_n003x = n5440_o; // (signal)
  /* vlm5030_gl.vhd:958:33  */
  assign start_block_n004x = n5443_o; // (signal)
  /* vlm5030_gl.vhd:958:40  */
  assign start_block_n005x = n5452_o; // (signal)
  /* vlm5030_gl.vhd:958:47  */
  assign start_block_n006x = n5453_o; // (signal)
  /* vlm5030_gl.vhd:959:12  */
  assign start_block_n007x = n5459_o; // (signal)
  /* vlm5030_gl.vhd:959:19  */
  assign start_block_n008x = n5463_o; // (signal)
  /* vlm5030_gl.vhd:959:26  */
  assign start_block_n009x = n5470_o; // (signal)
  /* vlm5030_gl.vhd:959:33  */
  assign start_block_n014x = n5530_o; // (signal)
  /* vlm5030_gl.vhd:959:40  */
  assign start_block_n015x = n5539_o; // (signal)
  /* vlm5030_gl.vhd:960:12  */
  assign start_block_n016x = n5548_o; // (signal)
  /* vlm5030_gl.vhd:960:19  */
  assign start_block_n017x = n5554_o; // (signal)
  /* vlm5030_gl.vhd:961:12  */
  assign start_block_n012x = n5526_o; // (signal)
  /* vlm5030_gl.vhd:963:12  */
  assign start_block_busy1q = n5748_q; // (signal)
  /* vlm5030_gl.vhd:964:12  */
  assign start_block_busy2q = n5750_q; // (signal)
  /* vlm5030_gl.vhd:965:12  */
  assign start_block_setbusy1 = n5632_o; // (signal)
  /* vlm5030_gl.vhd:968:16  */
  assign n5233_o = ~i_vcu;
  /* vlm5030_gl.vhd:969:16  */
  assign n5234_o = ~start_block_ffs1q;
  /* vlm5030_gl.vhd:971:17  */
  assign n5235_o = ~nvcufinal;
  assign n5243_o = clk2ena[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5245_o = clk2ena[2];
  /* vlm5030_gl.vhd:980:29  */
  assign n5247_o = start_block_startq[1:0];
  /* vlm5030_gl.vhd:980:42  */
  assign n5248_o = {n5247_o, starttst};
  /* vlm5030_gl.vhd:981:33  */
  assign n5249_o = ~(startrise & i_vcu);
  assign n5257_o = start_block_startq[1];
  /* vlm5030_gl.vhd:986:19  */
  assign n5258_o = ~n5257_o;
  assign n5259_o = start_block_startq[2];
  /* vlm5030_gl.vhd:986:32  */
  assign n5260_o = ~(n5258_o | n5259_o);
  /* vlm5030_gl.vhd:987:22  */
  assign n5261_o = ~start_block_startriseq;
  /* vlm5030_gl.vhd:990:22  */
  assign n5262_o = rstdel | start_block_n005x;
  assign n5270_o = clk2ena[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5272_o = clk2ena[2];
  /* vlm5030_gl.vhd:999:27  */
  assign n5274_o = start_block_ffs1nq & start_block_ffsloop;
  /* vlm5030_gl.vhd:999:55  */
  assign n5275_o = start_block_nvcu & startrise;
  /* vlm5030_gl.vhd:999:42  */
  assign n5276_o = ~(n5274_o | n5275_o);
  /* vlm5030_gl.vhd:1000:27  */
  assign n5277_o = start_block_ffs2nq & start_block_ffsloop;
  /* vlm5030_gl.vhd:1000:55  */
  assign n5278_o = i_vcu & startrise;
  /* vlm5030_gl.vhd:1000:42  */
  assign n5279_o = ~(n5277_o | n5278_o);
  /* vlm5030_gl.vhd:1001:27  */
  assign n5280_o = ~(start_block_ffs4q | startrise);
  assign n5281_o = start_block_startq[1];
  /* vlm5030_gl.vhd:1001:56  */
  assign n5282_o = ~(n5281_o | start_block_ffs3nq);
  /* vlm5030_gl.vhd:1001:42  */
  assign n5283_o = ~(n5280_o | n5282_o);
  /* vlm5030_gl.vhd:1002:26  */
  assign n5284_o = ~(start_block_ffs5nq & start_block_ffsloop);
  assign n5304_o = clk2ena[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5306_o = clk2ena[2];
  /* vlm5030_gl.vhd:1012:15  */
  assign n5310_o = ~start_block_ffs1q;
  /* vlm5030_gl.vhd:1013:15  */
  assign n5311_o = ~start_block_ffs2q;
  /* vlm5030_gl.vhd:1014:15  */
  assign n5312_o = ~start_block_ffs3q;
  /* vlm5030_gl.vhd:1015:15  */
  assign n5313_o = ~start_block_ffs4q;
  /* vlm5030_gl.vhd:1016:15  */
  assign n5314_o = ~start_block_ffs5q;
  /* vlm5030_gl.vhd:1018:26  */
  assign n5315_o = ~start_block_ffs3q;
  /* vlm5030_gl.vhd:1018:22  */
  assign n5316_o = start_block_ffs1q | n5315_o;
  /* vlm5030_gl.vhd:1018:52  */
  assign n5317_o = fsromdo[6];
  /* vlm5030_gl.vhd:1018:41  */
  assign n5318_o = ~n5317_o;
  /* vlm5030_gl.vhd:1018:37  */
  assign n5319_o = n5316_o | n5318_o;
  assign n5327_o = clk2enb[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5329_o = clk2enb[2];
  /* clock_functions_pack.vhd:65:34  */
  assign n5330_o = n5329_o & start_block_vcufinal1q;
  /* vlm5030_gl.vhd:1028:23  */
  assign n5331_o = ~start_block_vcufinal1q;
  /* vlm5030_gl.vhd:1031:25  */
  assign n5332_o = ~start_block_vcufinal2q;
  /* vlm5030_gl.vhd:1037:21  */
  assign n5341_o = ~start_block_vcufinal1q;
  /* vlm5030_gl.vhd:1037:42  */
  assign n5342_o = ~start_block_vcufinal2q;
  /* vlm5030_gl.vhd:1037:37  */
  assign n5343_o = ~(n5341_o | n5342_o);
  /* vlm5030_gl.vhd:1038:20  */
  assign n5344_o = ~vcufinal12;
  /* vlm5030_gl.vhd:1039:46  */
  assign n5345_o = ~start_block_ffs4q;
  /* vlm5030_gl.vhd:1039:41  */
  assign n5346_o = ~(start_block_ffs1q | n5345_o);
  /* vlm5030_gl.vhd:1039:27  */
  assign n5347_o = ~(rstdel | n5346_o);
  /* vlm5030_gl.vhd:1041:32  */
  assign n5348_o = ~(start_block_ffs3q | start_block_ffs1q);
  /* vlm5030_gl.vhd:1041:21  */
  assign n5349_o = start_block_ffs2nq ^ n5348_o;
  /* vlm5030_gl.vhd:1043:63  */
  assign n5350_o = fsromdo[6];
  /* vlm5030_gl.vhd:1043:52  */
  assign n5351_o = ~n5350_o;
  /* vlm5030_gl.vhd:1043:48  */
  assign n5352_o = start_block_ffs2nq | n5351_o;
  /* vlm5030_gl.vhd:1043:68  */
  assign n5353_o = n5352_o | start_block_nvcufinal12;
  /* vlm5030_gl.vhd:1043:36  */
  assign n5354_o = start_block_ffs3q & n5353_o;
  /* vlm5030_gl.vhd:1043:26  */
  assign n5355_o = start_block_ffs1q | n5354_o;
  /* vlm5030_gl.vhd:1045:5  */
  vlm5030_delay_inv_2 start_block_xromdo7nqdel_b (
    .i_clk_base(n5356_o),
    .i_clk_val(n5357_o),
    .i_clk_rise(n5358_o),
    .i_clk_fall(n5359_o),
    .i_in(xromdo7q),
    .o_out(start_block_xromdo7nqdel_b_o_out));
  assign n5356_o = osc[0];
  assign n5357_o = osc[1];
  assign n5358_o = osc[2];
  assign n5359_o = osc[3];
  /* vlm5030_gl.vhd:1056:28  */
  assign n5361_o = xromdo7nq & start_block_xromdo7nqdel;
  /* vlm5030_gl.vhd:1056:58  */
  assign n5362_o = start_block_vcumode | start_block_startriseqvcu;
  /* vlm5030_gl.vhd:1056:45  */
  assign n5363_o = n5361_o & n5362_o;
  /* vlm5030_gl.vhd:1056:77  */
  assign n5364_o = ~(n5363_o | start_block_ffs4nq);
  /* vlm5030_gl.vhd:1058:42  */
  assign n5365_o = fsromdo[7];
  /* vlm5030_gl.vhd:1058:46  */
  assign n5366_o = n5365_o & start_block_ffs3q;
  /* vlm5030_gl.vhd:1058:56  */
  assign n5367_o = n5366_o & vcufinal12;
  /* vlm5030_gl.vhd:1058:31  */
  assign n5368_o = start_block_startriseqvcu | n5367_o;
  /* vlm5030_gl.vhd:1061:23  */
  assign n5369_o = rstdel | startrise;
  assign n5377_o = c2d0[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5379_o = c2d0[2];
  /* vlm5030_gl.vhd:1068:49  */
  assign n5381_o = xromdo[7];
  /* vlm5030_gl.vhd:1068:39  */
  assign n5382_o = start_block_pmsff3nq & n5381_o;
  /* vlm5030_gl.vhd:1068:25  */
  assign n5383_o = ~(start_block_n008x | n5382_o);
  /* vlm5030_gl.vhd:1071:16  */
  assign n5388_o = ~start_block_msff1q;
  assign n5396_o = c2d6[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5398_o = c2d6[2];
  /* vlm5030_gl.vhd:1078:38  */
  assign n5400_o = xromdo[1];
  /* vlm5030_gl.vhd:1078:42  */
  assign n5401_o = n5400_o & start_block_n007x;
  /* vlm5030_gl.vhd:1078:52  */
  assign n5402_o = n5401_o & start_block_pmsff3nq;
  /* vlm5030_gl.vhd:1078:27  */
  assign n5403_o = ~(start_block_msff2nq | n5402_o);
  /* vlm5030_gl.vhd:1081:16  */
  assign n5408_o = ~start_block_msff2q;
  assign n5416_o = c2d6[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5418_o = c2d6[2];
  /* vlm5030_gl.vhd:1086:37  */
  assign n5420_o = xromdo[0];
  /* vlm5030_gl.vhd:1086:27  */
  assign n5421_o = start_block_n007x & n5420_o;
  /* vlm5030_gl.vhd:1086:56  */
  assign n5422_o = start_block_pmsff3nq & start_block_msff1q;
  /* vlm5030_gl.vhd:1086:42  */
  assign n5423_o = ~(n5421_o | n5422_o);
  /* vlm5030_gl.vhd:1089:17  */
  assign n5426_o = ~start_block_pmsff3q;
  /* vlm5030_gl.vhd:1092:31  */
  assign n5427_o = fsromdo[7];
  /* vlm5030_gl.vhd:1092:20  */
  assign n5428_o = ~n5427_o;
  /* vlm5030_gl.vhd:1092:36  */
  assign n5429_o = n5428_o | start_block_nvcufinal12;
  /* vlm5030_gl.vhd:1092:51  */
  assign n5430_o = n5429_o | start_block_ffs2nq;
  /* vlm5030_gl.vhd:1092:61  */
  assign n5431_o = n5430_o | start_block_ffs3nq;
  /* vlm5030_gl.vhd:1092:14  */
  assign n5432_o = ~n5431_o;
  /* vlm5030_gl.vhd:1093:21  */
  assign n5433_o = dq[0];
  /* vlm5030_gl.vhd:1093:25  */
  assign n5434_o = n5433_o | start_block_vcufinal2q;
  /* vlm5030_gl.vhd:1093:39  */
  assign n5435_o = n5434_o | start_block_vcufinal1q;
  /* vlm5030_gl.vhd:1093:14  */
  assign n5436_o = ~n5435_o;
  /* vlm5030_gl.vhd:1094:30  */
  assign n5437_o = dq[1];
  /* vlm5030_gl.vhd:1094:25  */
  assign n5438_o = start_block_n002x | n5437_o;
  /* vlm5030_gl.vhd:1094:34  */
  assign n5439_o = n5438_o | start_block_n004x;
  /* vlm5030_gl.vhd:1094:14  */
  assign n5440_o = ~n5439_o;
  /* vlm5030_gl.vhd:1095:36  */
  assign n5441_o = dq[0];
  /* vlm5030_gl.vhd:1095:30  */
  assign n5442_o = ~n5441_o;
  /* vlm5030_gl.vhd:1095:25  */
  assign n5443_o = ~(start_block_vcufinal1q | n5442_o);
  /* vlm5030_gl.vhd:1096:26  */
  assign n5445_o = start_block_msff2q | start_block_n006x;
  /* clock_functions_pack.vhd:147:24  */
  assign n5450_o = nc2d6[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n5451_o = n5445_o | n5450_o;
  /* vlm5030_gl.vhd:1096:14  */
  assign n5452_o = ~n5451_o;
  /* vlm5030_gl.vhd:1097:20  */
  assign n5453_o = ~(start_block_n009x & cntdn0);
  /* vlm5030_gl.vhd:1098:25  */
  assign n5454_o = start_block_n003x | start_block_ffs5nq;
  /* vlm5030_gl.vhd:1098:46  */
  assign n5455_o = fsromdo[13];
  /* vlm5030_gl.vhd:1098:62  */
  assign n5456_o = dinalq[7];
  /* vlm5030_gl.vhd:1098:51  */
  assign n5457_o = ~(n5455_o & n5456_o);
  /* vlm5030_gl.vhd:1098:35  */
  assign n5458_o = n5454_o | n5457_o;
  /* vlm5030_gl.vhd:1098:14  */
  assign n5459_o = ~n5458_o;
  /* vlm5030_gl.vhd:1099:26  */
  assign n5460_o = start_block_msff1q | rstdel;
  /* vlm5030_gl.vhd:1099:40  */
  assign n5461_o = ~start_block_n006x;
  /* vlm5030_gl.vhd:1099:36  */
  assign n5462_o = n5460_o | n5461_o;
  /* vlm5030_gl.vhd:1099:14  */
  assign n5463_o = ~n5462_o;
  /* vlm5030_gl.vhd:1100:46  */
  assign n5464_o = fsromdo[6];
  /* vlm5030_gl.vhd:1100:35  */
  assign n5465_o = ~n5464_o;
  /* vlm5030_gl.vhd:1100:31  */
  assign n5466_o = start_block_nvcufinal12 | n5465_o;
  /* vlm5030_gl.vhd:1100:65  */
  assign n5467_o = xromdo[7];
  /* vlm5030_gl.vhd:1100:55  */
  assign n5468_o = ~n5467_o;
  /* vlm5030_gl.vhd:1100:51  */
  assign n5469_o = n5466_o | n5468_o;
  /* vlm5030_gl.vhd:1100:14  */
  assign n5470_o = ~n5469_o;
  /* clock_functions_pack.vhd:139:26  */
  assign n5479_o = nc2d10[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n5480_o = nc2d10[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n5481_o = n5480_o | start_block_n003x;
  /* clock_functions_pack.vhd:141:26  */
  assign n5482_o = nc2d10[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n5483_o = ~start_block_n003x;
  /* clock_functions_pack.vhd:141:31  */
  assign n5484_o = n5482_o & n5483_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n5485_o = nc2d10[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n5486_o = ~start_block_n003x;
  /* clock_functions_pack.vhd:142:31  */
  assign n5487_o = n5485_o & n5486_o;
  assign n5488_o = {n5487_o, n5484_o, n5481_o, n5479_o};
  /* clock_functions_pack.vhd:139:26  */
  assign n5493_o = n5488_o[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n5494_o = n5488_o[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n5495_o = n5494_o | fsromevalout;
  /* clock_functions_pack.vhd:141:26  */
  assign n5496_o = n5488_o[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n5497_o = ~fsromevalout;
  /* clock_functions_pack.vhd:141:31  */
  assign n5498_o = n5496_o & n5497_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n5499_o = n5488_o[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n5500_o = ~fsromevalout;
  /* clock_functions_pack.vhd:142:31  */
  assign n5501_o = n5499_o & n5500_o;
  assign n5502_o = {n5501_o, n5498_o, n5495_o, n5493_o};
  /* clock_functions_pack.vhd:139:26  */
  assign n5507_o = n5502_o[0];
  /* clock_functions_pack.vhd:140:26  */
  assign n5508_o = n5502_o[1];
  /* clock_functions_pack.vhd:140:30  */
  assign n5509_o = n5508_o | start_block_ffs5nq;
  /* clock_functions_pack.vhd:141:26  */
  assign n5510_o = n5502_o[2];
  /* clock_functions_pack.vhd:141:35  */
  assign n5511_o = ~start_block_ffs5nq;
  /* clock_functions_pack.vhd:141:31  */
  assign n5512_o = n5510_o & n5511_o;
  /* clock_functions_pack.vhd:142:26  */
  assign n5513_o = n5502_o[3];
  /* clock_functions_pack.vhd:142:35  */
  assign n5514_o = ~start_block_ffs5nq;
  /* clock_functions_pack.vhd:142:31  */
  assign n5515_o = n5513_o & n5514_o;
  assign n5516_o = {n5515_o, n5512_o, n5509_o, n5507_o};
  /* clock_functions_pack.vhd:75:25  */
  assign n5521_o = n5516_o[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n5522_o = n5516_o[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n5523_o = ~n5522_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n5524_o = n5516_o[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n5525_o = n5516_o[2];
  assign n5526_o = {n5525_o, n5524_o, n5523_o, n5521_o};
  /* vlm5030_gl.vhd:1102:35  */
  assign n5527_o = start_block_n003x | start_block_ffs5nq;
  /* vlm5030_gl.vhd:1102:45  */
  assign n5528_o = n5527_o | fsromnorhigh;
  /* vlm5030_gl.vhd:1102:24  */
  assign n5529_o = ~n5528_o;
  /* vlm5030_gl.vhd:1102:20  */
  assign n5530_o = ~(start_block_n001x | n5529_o);
  /* vlm5030_gl.vhd:1103:21  */
  assign n5531_o = dq[1];
  /* vlm5030_gl.vhd:1103:25  */
  assign n5532_o = n5531_o | start_block_n004x;
  /* vlm5030_gl.vhd:1103:59  */
  assign n5533_o = ~start_block_vcufinal1q;
  /* vlm5030_gl.vhd:1103:55  */
  assign n5534_o = start_block_vcufinal2q | n5533_o;
  /* vlm5030_gl.vhd:1103:80  */
  assign n5535_o = dq[0];
  /* vlm5030_gl.vhd:1103:75  */
  assign n5536_o = n5534_o | n5535_o;
  /* vlm5030_gl.vhd:1103:38  */
  assign n5537_o = ~n5536_o;
  /* vlm5030_gl.vhd:1103:34  */
  assign n5538_o = n5532_o | n5537_o;
  /* vlm5030_gl.vhd:1103:14  */
  assign n5539_o = ~n5538_o;
  /* vlm5030_gl.vhd:1104:26  */
  assign n5540_o = fsromdo[6];
  /* vlm5030_gl.vhd:1104:15  */
  assign n5541_o = ~n5540_o;
  /* vlm5030_gl.vhd:1104:43  */
  assign n5542_o = dq[1];
  /* vlm5030_gl.vhd:1104:47  */
  assign n5543_o = n5542_o | start_block_n017x;
  /* vlm5030_gl.vhd:1104:62  */
  assign n5544_o = dq[0];
  /* vlm5030_gl.vhd:1104:66  */
  assign n5545_o = n5544_o & start_block_vcufinal1q;
  /* vlm5030_gl.vhd:1104:56  */
  assign n5546_o = n5543_o | n5545_o;
  /* vlm5030_gl.vhd:1104:36  */
  assign n5547_o = ~n5546_o;
  /* vlm5030_gl.vhd:1104:31  */
  assign n5548_o = ~(n5541_o | n5547_o);
  /* vlm5030_gl.vhd:1105:21  */
  assign n5549_o = dq[0];
  /* vlm5030_gl.vhd:1105:29  */
  assign n5550_o = ~vcufinal12;
  /* vlm5030_gl.vhd:1105:25  */
  assign n5551_o = n5549_o | n5550_o;
  /* vlm5030_gl.vhd:1105:49  */
  assign n5552_o = ~start_block_vcufinal1q;
  /* vlm5030_gl.vhd:1105:45  */
  assign n5553_o = n5551_o | n5552_o;
  /* vlm5030_gl.vhd:1105:14  */
  assign n5554_o = ~n5553_o;
  /* vlm5030_gl.vhd:1107:28  */
  assign n5555_o = start_block_msff1nq & start_block_n009x;
  /* vlm5030_gl.vhd:1107:43  */
  assign n5556_o = ~cntdn0;
  /* vlm5030_gl.vhd:1107:38  */
  assign n5557_o = n5555_o & n5556_o;
  /* vlm5030_gl.vhd:1107:15  */
  assign n5558_o = ~n5557_o;
  /* vlm5030_gl.vhd:1109:25  */
  assign n5559_o = xromdo[5];
  /* vlm5030_gl.vhd:1109:29  */
  assign n5560_o = ~(n5559_o & start_block_pmsff3nq);
  /* clock_functions_pack.vhd:93:26  */
  assign n5567_o = c2d0[0];
  /* clock_functions_pack.vhd:94:26  */
  assign n5568_o = c2d0[1];
  /* clock_functions_pack.vhd:94:30  */
  assign n5569_o = n5568_o & start_block_msff1nq;
  /* clock_functions_pack.vhd:95:26  */
  assign n5570_o = c2d0[2];
  /* clock_functions_pack.vhd:95:31  */
  assign n5571_o = n5570_o & start_block_msff1nq;
  /* clock_functions_pack.vhd:96:26  */
  assign n5572_o = c2d0[3];
  /* clock_functions_pack.vhd:96:31  */
  assign n5573_o = n5572_o & start_block_msff1nq;
  assign n5574_o = {n5573_o, n5571_o, n5569_o, n5567_o};
  /* vlm5030_gl.vhd:1110:56  */
  assign n5576_o = xromdo[5];
  /* vlm5030_gl.vhd:1110:60  */
  assign n5577_o = n5576_o & start_block_pmsff3nq;
  /* clock_functions_pack.vhd:93:26  */
  assign n5582_o = c2d6[0];
  /* clock_functions_pack.vhd:94:26  */
  assign n5583_o = c2d6[1];
  /* clock_functions_pack.vhd:94:30  */
  assign n5584_o = n5583_o & n5577_o;
  /* clock_functions_pack.vhd:95:26  */
  assign n5585_o = c2d6[2];
  /* clock_functions_pack.vhd:95:31  */
  assign n5586_o = n5585_o & n5577_o;
  /* clock_functions_pack.vhd:96:26  */
  assign n5587_o = c2d6[3];
  /* clock_functions_pack.vhd:96:31  */
  assign n5588_o = n5587_o & n5577_o;
  assign n5589_o = {n5588_o, n5586_o, n5584_o, n5582_o};
  /* clock_functions_pack.vhd:129:26  */
  assign n5594_o = n5574_o[0];
  /* clock_functions_pack.vhd:130:26  */
  assign n5595_o = n5574_o[1];
  /* clock_functions_pack.vhd:130:38  */
  assign n5596_o = n5589_o[1];
  /* clock_functions_pack.vhd:130:30  */
  assign n5597_o = n5595_o | n5596_o;
  /* clock_functions_pack.vhd:131:27  */
  assign n5598_o = n5574_o[2];
  /* clock_functions_pack.vhd:131:45  */
  assign n5599_o = n5589_o[1];
  /* clock_functions_pack.vhd:131:36  */
  assign n5600_o = ~n5599_o;
  /* clock_functions_pack.vhd:131:32  */
  assign n5601_o = n5598_o & n5600_o;
  /* clock_functions_pack.vhd:132:27  */
  assign n5602_o = n5589_o[2];
  /* clock_functions_pack.vhd:132:45  */
  assign n5603_o = n5574_o[1];
  /* clock_functions_pack.vhd:132:36  */
  assign n5604_o = ~n5603_o;
  /* clock_functions_pack.vhd:132:32  */
  assign n5605_o = n5602_o & n5604_o;
  /* clock_functions_pack.vhd:131:50  */
  assign n5606_o = n5601_o | n5605_o;
  /* clock_functions_pack.vhd:133:27  */
  assign n5607_o = n5574_o[3];
  /* clock_functions_pack.vhd:133:45  */
  assign n5608_o = n5589_o[1];
  /* clock_functions_pack.vhd:133:36  */
  assign n5609_o = ~n5608_o;
  /* clock_functions_pack.vhd:133:32  */
  assign n5610_o = n5607_o & n5609_o;
  /* clock_functions_pack.vhd:133:62  */
  assign n5611_o = n5589_o[2];
  /* clock_functions_pack.vhd:133:53  */
  assign n5612_o = ~n5611_o;
  /* clock_functions_pack.vhd:133:49  */
  assign n5613_o = n5610_o & n5612_o;
  /* clock_functions_pack.vhd:134:27  */
  assign n5614_o = n5589_o[3];
  /* clock_functions_pack.vhd:134:45  */
  assign n5615_o = n5574_o[1];
  /* clock_functions_pack.vhd:134:36  */
  assign n5616_o = ~n5615_o;
  /* clock_functions_pack.vhd:134:32  */
  assign n5617_o = n5614_o & n5616_o;
  /* clock_functions_pack.vhd:134:62  */
  assign n5618_o = n5574_o[2];
  /* clock_functions_pack.vhd:134:53  */
  assign n5619_o = ~n5618_o;
  /* clock_functions_pack.vhd:134:49  */
  assign n5620_o = n5617_o & n5619_o;
  /* clock_functions_pack.vhd:133:68  */
  assign n5621_o = n5613_o | n5620_o;
  assign n5622_o = {n5621_o, n5606_o, n5597_o, n5594_o};
  /* clock_functions_pack.vhd:147:24  */
  assign n5628_o = start_block_n012x[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n5629_o = start_block_msff1nq | n5628_o;
  /* vlm5030_gl.vhd:1114:20  */
  assign n5630_o = ~(start_block_n014x | start_block_msff1nq);
  assign n5631_o = start_block_startq[1];
  /* vlm5030_gl.vhd:1117:25  */
  assign n5632_o = ~(n5631_o | start_block_startriseqvcu);
  assign n5640_o = clk2ctrl[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5642_o = clk2ctrl[2];
  /* vlm5030_gl.vhd:1123:38  */
  assign n5644_o = ~start_block_busy1q;
  /* vlm5030_gl.vhd:1123:33  */
  assign n5645_o = ~(start_block_startriseqvcu | n5644_o);
  assign n5657_o = clk2ctrl[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5659_o = clk2ctrl[2];
  /* vlm5030_gl.vhd:1132:32  */
  assign n5661_o = ~start_block_busy2q;
  /* vlm5030_gl.vhd:1132:27  */
  assign n5662_o = ~(start_block_vcumode | n5661_o);
  /* vlm5030_gl.vhd:1136:14  */
  assign n5667_o = ~start_block_busy1q;
  /* vlm5030_gl.vhd:1136:31  */
  assign n5668_o = ~start_block_busy2q;
  /* vlm5030_gl.vhd:1136:26  */
  assign n5669_o = ~(n5667_o | n5668_o);
  /* vlm5030_gl.vhd:1138:22  */
  assign n5670_o = start_block_ffs4q | i_start;
  /* vlm5030_gl.vhd:1138:33  */
  assign n5671_o = n5670_o | xromdo7nq;
  /* vlm5030_gl.vhd:1138:11  */
  assign n5672_o = ~n5671_o;
  /* vlm5030_gl.vhd:1140:37  */
  assign n5674_o = fsromevalout | start_block_n003x;
  /* clock_functions_pack.vhd:147:24  */
  assign n5679_o = nc2d6[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n5680_o = n5674_o | n5679_o;
  /* vlm5030_gl.vhd:1140:19  */
  assign n5681_o = ~n5680_o;
  /* vlm5030_gl.vhd:1142:38  */
  assign n5682_o = dq[1];
  /* vlm5030_gl.vhd:1142:33  */
  assign n5683_o = start_block_vcufinal2q | n5682_o;
  /* vlm5030_gl.vhd:1142:47  */
  assign n5684_o = dq[0];
  /* vlm5030_gl.vhd:1142:42  */
  assign n5685_o = n5683_o | n5684_o;
  /* vlm5030_gl.vhd:1142:17  */
  assign n5686_o = ~n5685_o;
  /* vlm5030_gl.vhd:1144:44  */
  assign n5687_o = fsromdo[6];
  /* vlm5030_gl.vhd:1144:33  */
  assign n5688_o = ~n5687_o;
  /* vlm5030_gl.vhd:1144:29  */
  assign n5689_o = start_block_n015x | n5688_o;
  /* vlm5030_gl.vhd:1144:63  */
  assign n5690_o = xromdo[11];
  /* vlm5030_gl.vhd:1144:53  */
  assign n5691_o = ~n5690_o;
  /* vlm5030_gl.vhd:1144:49  */
  assign n5692_o = n5689_o | n5691_o;
  /* vlm5030_gl.vhd:1144:18  */
  assign n5693_o = ~n5692_o;
  /* vlm5030_gl.vhd:1146:43  */
  assign n5695_o = ~(tstend2id | start_block_ffs5nq);
  /* vlm5030_gl.vhd:1146:28  */
  assign n5696_o = start_block_n016x & n5695_o;
  /* vlm5030_gl.vhd:1146:17  */
  assign n5697_o = ~n5696_o;
  /* clock_functions_pack.vhd:170:25  */
  assign n5702_o = nc2d8[1];
  /* clock_functions_pack.vhd:170:16  */
  assign n5703_o = ~(n5697_o | n5702_o);
  /* vlm5030_gl.vhd:1150:29  */
  assign n5704_o = start_block_ffs5nq | tstend2id;
  /* clock_functions_pack.vhd:170:25  */
  assign n5711_o = nc2d8[1];
  /* clock_functions_pack.vhd:170:16  */
  assign n5712_o = ~(start_block_n016x | n5711_o);
  /* clock_functions_pack.vhd:170:25  */
  assign n5717_o = c2d4[1];
  /* clock_functions_pack.vhd:170:16  */
  assign n5718_o = ~(n5712_o | n5717_o);
  /* vlm5030_gl.vhd:1150:42  */
  assign n5719_o = n5704_o | n5718_o;
  /* vlm5030_gl.vhd:1150:17  */
  assign n5720_o = ~n5719_o;
  /* vlm5030_gl.vhd:979:7  */
  assign n5721_o = n5245_o ? n5248_o : start_block_startq;
  /* vlm5030_gl.vhd:979:7  */
  always @(posedge n5243_o or posedge rstdel)
    if (rstdel)
      n5722_q <= 3'b000;
    else
      n5722_q <= n5721_o;
  /* vlm5030_gl.vhd:979:7  */
  assign n5723_o = n5245_o ? n5249_o : start_block_startriseq;
  /* vlm5030_gl.vhd:979:7  */
  always @(posedge n5243_o or posedge rstdel)
    if (rstdel)
      n5724_q <= 1'b1;
    else
      n5724_q <= n5723_o;
  /* vlm5030_gl.vhd:998:7  */
  assign n5725_o = n5272_o ? n5276_o : start_block_ffs1q;
  /* vlm5030_gl.vhd:998:7  */
  always @(posedge n5270_o or posedge start_block_ffsset)
    if (start_block_ffsset)
      n5726_q <= 1'b1;
    else
      n5726_q <= n5725_o;
  /* vlm5030_gl.vhd:991:5  */
  assign n5727_o = ~start_block_ffsset;
  /* vlm5030_gl.vhd:991:5  */
  assign n5728_o = n5272_o & n5727_o;
  /* vlm5030_gl.vhd:998:7  */
  assign n5729_o = n5728_o ? n5279_o : start_block_ffs2q;
  /* vlm5030_gl.vhd:998:7  */
  always @(posedge n5270_o)
    n5730_q <= n5729_o;
  initial
    n5730_q = 1'b1;
  /* vlm5030_gl.vhd:1008:7  */
  assign n5731_o = n5306_o ? start_block_ffs1nq : start_block_ffs3q;
  /* vlm5030_gl.vhd:1008:7  */
  always @(posedge n5304_o)
    n5732_q <= n5731_o;
  initial
    n5732_q = 1'b1;
  /* vlm5030_gl.vhd:998:7  */
  assign n5733_o = n5272_o ? n5283_o : start_block_ffs4q;
  /* vlm5030_gl.vhd:998:7  */
  always @(posedge n5270_o or posedge start_block_ffsset)
    if (start_block_ffsset)
      n5734_q <= 1'b1;
    else
      n5734_q <= n5733_o;
  /* vlm5030_gl.vhd:998:7  */
  assign n5735_o = n5272_o ? n5284_o : start_block_ffs5q;
  /* vlm5030_gl.vhd:998:7  */
  always @(posedge n5270_o or posedge start_block_ffsset)
    if (start_block_ffsset)
      n5736_q <= 1'b0;
    else
      n5736_q <= n5735_o;
  /* vlm5030_gl.vhd:1027:7  */
  assign n5737_o = n5329_o ? n5331_o : start_block_vcufinal1q;
  /* vlm5030_gl.vhd:1027:7  */
  always @(posedge n5327_o or posedge start_block_vcufinal)
    if (start_block_vcufinal)
      n5738_q <= 1'b1;
    else
      n5738_q <= n5737_o;
  /* vlm5030_gl.vhd:1027:7  */
  assign n5739_o = n5330_o ? n5332_o : start_block_vcufinal2q;
  /* vlm5030_gl.vhd:1027:7  */
  always @(posedge n5327_o or posedge start_block_vcufinal)
    if (start_block_vcufinal)
      n5740_q <= 1'b1;
    else
      n5740_q <= n5739_o;
  /* vlm5030_gl.vhd:1067:7  */
  assign n5741_o = n5379_o ? n5383_o : start_block_msff1q;
  /* vlm5030_gl.vhd:1067:7  */
  always @(posedge n5377_o or posedge start_block_msffset)
    if (start_block_msffset)
      n5742_q <= 1'b1;
    else
      n5742_q <= n5741_o;
  /* vlm5030_gl.vhd:1077:7  */
  assign n5743_o = n5398_o ? n5403_o : start_block_msff2q;
  /* vlm5030_gl.vhd:1077:7  */
  always @(posedge n5396_o or posedge start_block_msffset)
    if (start_block_msffset)
      n5744_q <= 1'b1;
    else
      n5744_q <= n5743_o;
  /* vlm5030_gl.vhd:1085:7  */
  assign n5745_o = n5418_o ? n5423_o : start_block_pmsff3q;
  /* vlm5030_gl.vhd:1085:7  */
  always @(posedge n5416_o)
    n5746_q <= n5745_o;
  initial
    n5746_q = 1'b0;
  /* vlm5030_gl.vhd:1122:7  */
  assign n5747_o = n5642_o ? n5645_o : start_block_busy1q;
  /* vlm5030_gl.vhd:1122:7  */
  always @(posedge n5640_o or posedge start_block_setbusy1)
    if (start_block_setbusy1)
      n5748_q <= 1'b1;
    else
      n5748_q <= n5747_o;
  /* vlm5030_gl.vhd:1131:7  */
  assign n5749_o = n5659_o ? n5662_o : start_block_busy2q;
  /* vlm5030_gl.vhd:1131:7  */
  always @(posedge n5657_o or posedge start_block_ffsset)
    if (start_block_ffsset)
      n5750_q <= 1'b1;
    else
      n5750_q <= n5749_o;
  /* vlm5030_gl.vhd:1160:12  */
  assign krom_block_ka = n5751_o; // (signal)
  /* vlm5030_gl.vhd:1164:14  */
  assign krom_block_agen_block_nfsrdo6 = n5831_o; // (signal)
  /* vlm5030_gl.vhd:1165:14  */
  assign krom_block_agen_block_ksaq = n5863_q; // (signal)
  /* vlm5030_gl.vhd:1168:20  */
  assign n5751_o = dinalq[7:3];
  /* vlm5030_gl.vhd:1171:18  */
  always @*
    krom_block_agen_block_n5752_toggle = n5829_q; // (isignal)
  initial
    krom_block_agen_block_n5752_toggle = 5'bX;
  /* vlm5030_gl.vhd:1173:19  */
  assign n5755_o = fsromdo[6];
  assign n5761_o = clkksa[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n5763_o = clkksa[2];
  assign n5766_o = krom_block_agen_block_n5752_toggle[4:1];
  assign n5767_o = {n5766_o, 1'b1};
  /* vlm5030_gl.vhd:1179:22  */
  assign n5768_o = n5767_o[0];
  /* vlm5030_gl.vhd:1180:36  */
  assign n5769_o = krom_block_agen_block_ksaq[0];
  /* vlm5030_gl.vhd:1180:28  */
  assign n5770_o = ~n5769_o;
  assign n5771_o = krom_block_agen_block_ksaq[0];
  /* vlm5030_gl.vhd:1179:13  */
  assign n5772_o = n5768_o ? n5770_o : n5771_o;
  /* vlm5030_gl.vhd:1183:34  */
  assign n5773_o = krom_block_agen_block_ksaq[0];
  assign n5774_o = krom_block_agen_block_n5752_toggle[4:1];
  assign n5775_o = {n5774_o, 1'b1};
  /* vlm5030_gl.vhd:1183:55  */
  assign n5776_o = n5775_o[0];
  /* vlm5030_gl.vhd:1183:45  */
  assign n5777_o = ~n5776_o;
  /* vlm5030_gl.vhd:1183:40  */
  assign n5778_o = ~(n5773_o | n5777_o);
  assign n5779_o = krom_block_agen_block_n5752_toggle[4:2];
  assign n5780_o = {n5779_o, n5778_o, 1'b1};
  /* vlm5030_gl.vhd:1179:22  */
  assign n5781_o = n5780_o[1];
  /* vlm5030_gl.vhd:1180:36  */
  assign n5782_o = krom_block_agen_block_ksaq[1];
  /* vlm5030_gl.vhd:1180:28  */
  assign n5783_o = ~n5782_o;
  assign n5784_o = krom_block_agen_block_ksaq[1];
  /* vlm5030_gl.vhd:1179:13  */
  assign n5785_o = n5781_o ? n5783_o : n5784_o;
  /* vlm5030_gl.vhd:1183:34  */
  assign n5786_o = krom_block_agen_block_ksaq[1];
  assign n5787_o = krom_block_agen_block_n5752_toggle[4:2];
  assign n5788_o = {n5787_o, n5778_o, 1'b1};
  /* vlm5030_gl.vhd:1183:55  */
  assign n5789_o = n5788_o[1];
  /* vlm5030_gl.vhd:1183:45  */
  assign n5790_o = ~n5789_o;
  /* vlm5030_gl.vhd:1183:40  */
  assign n5791_o = ~(n5786_o | n5790_o);
  assign n5792_o = krom_block_agen_block_n5752_toggle[4:3];
  assign n5793_o = {n5792_o, n5791_o, n5778_o, 1'b1};
  /* vlm5030_gl.vhd:1179:22  */
  assign n5794_o = n5793_o[2];
  /* vlm5030_gl.vhd:1180:36  */
  assign n5795_o = krom_block_agen_block_ksaq[2];
  /* vlm5030_gl.vhd:1180:28  */
  assign n5796_o = ~n5795_o;
  assign n5797_o = krom_block_agen_block_ksaq[2];
  /* vlm5030_gl.vhd:1179:13  */
  assign n5798_o = n5794_o ? n5796_o : n5797_o;
  /* vlm5030_gl.vhd:1183:34  */
  assign n5799_o = krom_block_agen_block_ksaq[2];
  assign n5800_o = krom_block_agen_block_n5752_toggle[4:3];
  assign n5801_o = {n5800_o, n5791_o, n5778_o, 1'b1};
  /* vlm5030_gl.vhd:1183:55  */
  assign n5802_o = n5801_o[2];
  /* vlm5030_gl.vhd:1183:45  */
  assign n5803_o = ~n5802_o;
  /* vlm5030_gl.vhd:1183:40  */
  assign n5804_o = ~(n5799_o | n5803_o);
  assign n5805_o = krom_block_agen_block_n5752_toggle[4];
  assign n5806_o = {n5805_o, n5804_o, n5791_o, n5778_o, 1'b1};
  /* vlm5030_gl.vhd:1179:22  */
  assign n5807_o = n5806_o[3];
  /* vlm5030_gl.vhd:1180:36  */
  assign n5808_o = krom_block_agen_block_ksaq[3];
  /* vlm5030_gl.vhd:1180:28  */
  assign n5809_o = ~n5808_o;
  assign n5810_o = krom_block_agen_block_ksaq[3];
  /* vlm5030_gl.vhd:1179:13  */
  assign n5811_o = n5807_o ? n5809_o : n5810_o;
  /* vlm5030_gl.vhd:1183:34  */
  assign n5812_o = krom_block_agen_block_ksaq[3];
  assign n5813_o = krom_block_agen_block_n5752_toggle[4];
  assign n5814_o = {n5813_o, n5804_o, n5791_o, n5778_o, 1'b1};
  /* vlm5030_gl.vhd:1183:55  */
  assign n5815_o = n5814_o[3];
  /* vlm5030_gl.vhd:1183:45  */
  assign n5816_o = ~n5815_o;
  /* vlm5030_gl.vhd:1183:40  */
  assign n5817_o = ~(n5812_o | n5816_o);
  assign n5818_o = {n5811_o, n5798_o, n5785_o, n5772_o};
  assign n5820_o = {n5817_o, n5804_o, n5791_o, n5778_o, 1'b1};
  /* vlm5030_gl.vhd:1170:7  */
  assign n5826_o = ~n5755_o;
  /* vlm5030_gl.vhd:1170:7  */
  assign n5827_o = n5763_o & n5826_o;
  /* vlm5030_gl.vhd:1176:9  */
  assign n5828_o = n5827_o ? n5820_o : krom_block_agen_block_n5752_toggle;
  /* vlm5030_gl.vhd:1176:9  */
  always @(posedge n5761_o)
    n5829_q <= n5828_o;
  /* vlm5030_gl.vhd:1189:29  */
  assign n5830_o = fsromdo[6];
  /* vlm5030_gl.vhd:1189:18  */
  assign n5831_o = ~n5830_o;
  /* vlm5030_gl.vhd:1192:24  */
  assign n5832_o = krom_block_agen_block_ksaq[0];
  /* vlm5030_gl.vhd:1192:16  */
  assign n5833_o = ~n5832_o;
  /* vlm5030_gl.vhd:1192:29  */
  assign n5834_o = n5833_o & krom_block_agen_block_nfsrdo6;
  /* vlm5030_gl.vhd:1192:65  */
  assign n5835_o = yromdo[3];
  /* vlm5030_gl.vhd:1192:55  */
  assign n5836_o = ~(krom_block_agen_block_nfsrdo6 | n5835_o);
  /* vlm5030_gl.vhd:1192:42  */
  assign n5837_o = ~(n5834_o | n5836_o);
  /* vlm5030_gl.vhd:1193:24  */
  assign n5838_o = krom_block_agen_block_ksaq[1];
  /* vlm5030_gl.vhd:1193:16  */
  assign n5839_o = ~n5838_o;
  /* vlm5030_gl.vhd:1193:29  */
  assign n5840_o = n5839_o & krom_block_agen_block_nfsrdo6;
  /* vlm5030_gl.vhd:1193:65  */
  assign n5841_o = yromdo[2];
  /* vlm5030_gl.vhd:1193:55  */
  assign n5842_o = ~(krom_block_agen_block_nfsrdo6 | n5841_o);
  /* vlm5030_gl.vhd:1193:42  */
  assign n5843_o = ~(n5840_o | n5842_o);
  /* vlm5030_gl.vhd:1194:24  */
  assign n5844_o = krom_block_agen_block_ksaq[2];
  /* vlm5030_gl.vhd:1194:16  */
  assign n5845_o = ~n5844_o;
  /* vlm5030_gl.vhd:1194:29  */
  assign n5846_o = n5845_o & krom_block_agen_block_nfsrdo6;
  /* vlm5030_gl.vhd:1194:65  */
  assign n5847_o = yromdo[1];
  /* vlm5030_gl.vhd:1194:55  */
  assign n5848_o = ~(krom_block_agen_block_nfsrdo6 | n5847_o);
  /* vlm5030_gl.vhd:1194:42  */
  assign n5849_o = ~(n5846_o | n5848_o);
  /* vlm5030_gl.vhd:1195:24  */
  assign n5850_o = krom_block_agen_block_ksaq[3];
  /* vlm5030_gl.vhd:1195:16  */
  assign n5851_o = ~n5850_o;
  /* vlm5030_gl.vhd:1195:29  */
  assign n5852_o = n5851_o & krom_block_agen_block_nfsrdo6;
  /* vlm5030_gl.vhd:1195:54  */
  assign n5853_o = fsromdo[6];
  /* vlm5030_gl.vhd:1195:69  */
  assign n5854_o = yromdo[0];
  /* vlm5030_gl.vhd:1195:84  */
  assign n5855_o = xromdo[10];
  /* vlm5030_gl.vhd:1195:99  */
  assign n5856_o = xromdo[11];
  /* vlm5030_gl.vhd:1195:89  */
  assign n5857_o = ~(n5855_o | n5856_o);
  /* vlm5030_gl.vhd:1195:73  */
  assign n5858_o = n5854_o ^ n5857_o;
  /* vlm5030_gl.vhd:1195:58  */
  assign n5859_o = n5853_o & n5858_o;
  /* vlm5030_gl.vhd:1195:42  */
  assign n5860_o = ~(n5852_o | n5859_o);
  assign n5861_o = {n5860_o, n5849_o, n5843_o, n5837_o};
  /* vlm5030_gl.vhd:1176:9  */
  assign n5862_o = n5763_o ? n5818_o : krom_block_agen_block_ksaq;
  /* vlm5030_gl.vhd:1176:9  */
  always @(posedge n5761_o or posedge n5755_o)
    if (n5755_o)
      n5863_q <= 4'b1011;
    else
      n5863_q <= n5862_o;
  /* vlm5030_gl.vhd:1201:14  */
  assign krom_block_rom_block_kslice0 = n7308_o; // (signal)
  /* vlm5030_gl.vhd:1201:23  */
  assign krom_block_rom_block_kslice1 = n8742_o; // (signal)
  /* vlm5030_gl.vhd:1201:32  */
  assign krom_block_rom_block_kslice2 = n10176_o; // (signal)
  /* vlm5030_gl.vhd:1201:41  */
  assign krom_block_rom_block_kslice3 = n11184_o; // (signal)
  /* vlm5030_gl.vhd:1201:50  */
  assign krom_block_rom_block_kslice4 = n12192_o; // (signal)
  /* vlm5030_gl.vhd:1201:59  */
  assign krom_block_rom_block_kslice5 = n12210_o; // (signal)
  /* vlm5030_gl.vhd:1204:14  */
  assign krom_block_rom_block_wl = n20542_o; // (signal)
  /* vlm5030_gl.vhd:1205:14  */
  assign krom_block_rom_block_wl_slice = n12251_o; // (signal)
  /* vlm5030_gl.vhd:1208:14  */
  assign krom_block_rom_block_nkaodd = n12233_o; // (signal)
  /* vlm5030_gl.vhd:1210:14  */
  assign krom_block_rom_block_nksa0 = n12235_o; // (signal)
  /* vlm5030_gl.vhd:1211:14  */
  assign krom_block_rom_block_range_s0s1s2 = n12226_o; // (signal)
  /* vlm5030_gl.vhd:1211:28  */
  assign krom_block_rom_block_range_s3s4 = n12231_o; // (signal)
  /* vlm5030_gl.vhd:1213:14  */
  assign krom_block_rom_block_kout = n12693_o; // (signal)
  /* vlm5030_gl.vhd:1219:12  */
  assign n5868_o = 5'b11111 - krom_block_ka;
  /* vlm5030_pack.vhd:50:26  */
  assign n5886_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n5888_o = n5886_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5890_o = 1'b0 | n5888_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5892_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n5894_o = n5892_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5895_o = n5890_o | n5894_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5896_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n5898_o = n5896_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5899_o = n5895_o | n5898_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5900_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n5902_o = n5900_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5903_o = n5899_o | n5902_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5904_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n5906_o = n5904_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5907_o = n5903_o | n5906_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5908_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n5910_o = n5908_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5911_o = n5907_o | n5910_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5912_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n5914_o = n5912_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5915_o = n5911_o | n5914_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5916_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n5918_o = n5916_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5919_o = n5915_o | n5918_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5920_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n5922_o = n5920_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5923_o = n5919_o | n5922_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5924_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n5926_o = n5924_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5927_o = n5923_o | n5926_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5928_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n5930_o = n5928_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5931_o = n5927_o | n5930_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5932_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n5934_o = n5932_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5935_o = n5931_o | n5934_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5936_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n5938_o = n5936_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5939_o = n5935_o | n5938_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5940_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n5942_o = n5940_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5943_o = n5939_o | n5942_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5944_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n5946_o = n5944_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5947_o = n5943_o | n5946_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5948_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n5950_o = n5948_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5951_o = n5947_o | n5950_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5952_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n5954_o = n5952_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5955_o = n5951_o | n5954_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5956_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n5958_o = n5956_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5959_o = n5955_o | n5958_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5960_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n5962_o = n5960_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5963_o = n5959_o | n5962_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5964_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n5966_o = n5964_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5967_o = n5963_o | n5966_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5968_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n5970_o = n5968_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5971_o = n5967_o | n5970_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5972_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n5974_o = n5972_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5975_o = n5971_o | n5974_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5976_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n5978_o = n5976_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5979_o = n5975_o | n5978_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5980_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n5982_o = n5980_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5983_o = n5979_o | n5982_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5984_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n5986_o = n5984_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5987_o = n5983_o | n5986_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5988_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n5990_o = n5988_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n5991_o = n5987_o | n5990_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5992_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n5994_o = n5992_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5995_o = n5991_o | n5994_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n5996_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n5998_o = n5996_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n5999_o = n5995_o | n5998_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6000_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n6002_o = n6000_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6003_o = n5999_o | n6002_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6004_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n6006_o = n6004_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6007_o = n6003_o | n6006_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6008_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n6010_o = n6008_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6011_o = n6007_o | n6010_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6012_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n6014_o = n6012_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6015_o = n6011_o | n6014_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n6016_o = ~n6015_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n6017_o = ~n6016_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6029_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n6031_o = n6029_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6033_o = 1'b0 | n6031_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6035_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n6037_o = n6035_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6038_o = n6033_o | n6037_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6039_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n6041_o = n6039_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6042_o = n6038_o | n6041_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6043_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n6045_o = n6043_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6046_o = n6042_o | n6045_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6047_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n6049_o = n6047_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6050_o = n6046_o | n6049_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6051_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n6053_o = n6051_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6054_o = n6050_o | n6053_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6055_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n6057_o = n6055_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6058_o = n6054_o | n6057_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6059_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n6061_o = n6059_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6062_o = n6058_o | n6061_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6063_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n6065_o = n6063_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6066_o = n6062_o | n6065_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6067_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n6069_o = n6067_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6070_o = n6066_o | n6069_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6071_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n6073_o = n6071_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6074_o = n6070_o | n6073_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6075_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n6077_o = n6075_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6078_o = n6074_o | n6077_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6079_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n6081_o = n6079_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6082_o = n6078_o | n6081_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6083_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n6085_o = n6083_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6086_o = n6082_o | n6085_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6087_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n6089_o = n6087_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6090_o = n6086_o | n6089_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6091_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n6093_o = n6091_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6094_o = n6090_o | n6093_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6095_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n6097_o = n6095_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6098_o = n6094_o | n6097_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6099_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n6101_o = n6099_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6102_o = n6098_o | n6101_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6103_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n6105_o = n6103_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6106_o = n6102_o | n6105_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6107_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n6109_o = n6107_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6110_o = n6106_o | n6109_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6111_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n6113_o = n6111_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6114_o = n6110_o | n6113_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6115_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n6117_o = n6115_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6118_o = n6114_o | n6117_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6119_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n6121_o = n6119_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6122_o = n6118_o | n6121_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6123_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n6125_o = n6123_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6126_o = n6122_o | n6125_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6127_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n6129_o = n6127_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6130_o = n6126_o | n6129_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6131_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n6133_o = n6131_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6134_o = n6130_o | n6133_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6135_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n6137_o = n6135_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6138_o = n6134_o | n6137_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6139_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n6141_o = n6139_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6142_o = n6138_o | n6141_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6143_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n6145_o = n6143_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6146_o = n6142_o | n6145_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6147_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n6149_o = n6147_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6150_o = n6146_o | n6149_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6151_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n6153_o = n6151_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6154_o = n6150_o | n6153_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6155_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n6157_o = n6155_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6158_o = n6154_o | n6157_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n6159_o = ~n6158_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n6160_o = ~n6159_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6172_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n6174_o = n6172_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6176_o = 1'b0 | n6174_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6178_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n6180_o = n6178_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6181_o = n6176_o | n6180_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6182_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n6184_o = n6182_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6185_o = n6181_o | n6184_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6186_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n6188_o = n6186_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6189_o = n6185_o | n6188_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6190_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n6192_o = n6190_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6193_o = n6189_o | n6192_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6194_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n6196_o = n6194_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6197_o = n6193_o | n6196_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6198_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n6200_o = n6198_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6201_o = n6197_o | n6200_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6202_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n6204_o = n6202_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6205_o = n6201_o | n6204_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6206_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n6208_o = n6206_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6209_o = n6205_o | n6208_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6210_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n6212_o = n6210_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6213_o = n6209_o | n6212_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6214_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n6216_o = n6214_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6217_o = n6213_o | n6216_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6218_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n6220_o = n6218_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6221_o = n6217_o | n6220_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6222_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n6224_o = n6222_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6225_o = n6221_o | n6224_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6226_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n6228_o = n6226_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6229_o = n6225_o | n6228_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6230_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n6232_o = n6230_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6233_o = n6229_o | n6232_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6234_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n6236_o = n6234_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6237_o = n6233_o | n6236_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6238_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n6240_o = n6238_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6241_o = n6237_o | n6240_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6242_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n6244_o = n6242_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6245_o = n6241_o | n6244_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6246_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n6248_o = n6246_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6249_o = n6245_o | n6248_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6250_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n6252_o = n6250_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6253_o = n6249_o | n6252_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6254_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n6256_o = n6254_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6257_o = n6253_o | n6256_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6258_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n6260_o = n6258_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6261_o = n6257_o | n6260_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6262_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n6264_o = n6262_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6265_o = n6261_o | n6264_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6266_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n6268_o = n6266_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6269_o = n6265_o | n6268_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6270_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n6272_o = n6270_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6273_o = n6269_o | n6272_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6274_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n6276_o = n6274_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6277_o = n6273_o | n6276_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6278_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n6280_o = n6278_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6281_o = n6277_o | n6280_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6282_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n6284_o = n6282_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6285_o = n6281_o | n6284_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6286_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n6288_o = n6286_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6289_o = n6285_o | n6288_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6290_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n6292_o = n6290_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6293_o = n6289_o | n6292_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6294_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n6296_o = n6294_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6297_o = n6293_o | n6296_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6298_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n6300_o = n6298_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6301_o = n6297_o | n6300_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n6302_o = ~n6301_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n6303_o = ~n6302_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6315_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n6317_o = n6315_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6319_o = 1'b0 | n6317_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6321_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n6323_o = n6321_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6324_o = n6319_o | n6323_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6325_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n6327_o = n6325_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6328_o = n6324_o | n6327_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6329_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n6331_o = n6329_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6332_o = n6328_o | n6331_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6333_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n6335_o = n6333_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6336_o = n6332_o | n6335_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6337_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n6339_o = n6337_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6340_o = n6336_o | n6339_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6341_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n6343_o = n6341_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6344_o = n6340_o | n6343_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6345_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n6347_o = n6345_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6348_o = n6344_o | n6347_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6349_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n6351_o = n6349_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6352_o = n6348_o | n6351_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6353_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n6355_o = n6353_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6356_o = n6352_o | n6355_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6357_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n6359_o = n6357_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6360_o = n6356_o | n6359_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6361_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n6363_o = n6361_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6364_o = n6360_o | n6363_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6365_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n6367_o = n6365_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6368_o = n6364_o | n6367_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6369_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n6371_o = n6369_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6372_o = n6368_o | n6371_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6373_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n6375_o = n6373_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6376_o = n6372_o | n6375_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6377_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n6379_o = n6377_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6380_o = n6376_o | n6379_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6381_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n6383_o = n6381_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6384_o = n6380_o | n6383_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6385_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n6387_o = n6385_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6388_o = n6384_o | n6387_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6389_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n6391_o = n6389_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6392_o = n6388_o | n6391_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6393_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n6395_o = n6393_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6396_o = n6392_o | n6395_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6397_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n6399_o = n6397_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6400_o = n6396_o | n6399_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6401_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n6403_o = n6401_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6404_o = n6400_o | n6403_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6405_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n6407_o = n6405_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6408_o = n6404_o | n6407_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6409_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n6411_o = n6409_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6412_o = n6408_o | n6411_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6413_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n6415_o = n6413_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6416_o = n6412_o | n6415_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6417_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n6419_o = n6417_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6420_o = n6416_o | n6419_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6421_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n6423_o = n6421_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6424_o = n6420_o | n6423_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6425_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n6427_o = n6425_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6428_o = n6424_o | n6427_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6429_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n6431_o = n6429_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6432_o = n6428_o | n6431_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6433_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n6435_o = n6433_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6436_o = n6432_o | n6435_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6437_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n6439_o = n6437_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6440_o = n6436_o | n6439_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6441_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n6443_o = n6441_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6444_o = n6440_o | n6443_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n6445_o = ~n6444_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n6446_o = ~n6445_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6458_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n6460_o = n6458_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6462_o = 1'b0 | n6460_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6464_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n6466_o = n6464_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6467_o = n6462_o | n6466_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6468_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n6470_o = n6468_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6471_o = n6467_o | n6470_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6472_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n6474_o = n6472_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6475_o = n6471_o | n6474_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6476_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n6478_o = n6476_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6479_o = n6475_o | n6478_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6480_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n6482_o = n6480_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6483_o = n6479_o | n6482_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6484_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n6486_o = n6484_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6487_o = n6483_o | n6486_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6488_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n6490_o = n6488_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6491_o = n6487_o | n6490_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6492_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n6494_o = n6492_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6495_o = n6491_o | n6494_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6496_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n6498_o = n6496_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6499_o = n6495_o | n6498_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6500_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n6502_o = n6500_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6503_o = n6499_o | n6502_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6504_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n6506_o = n6504_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6507_o = n6503_o | n6506_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6508_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n6510_o = n6508_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6511_o = n6507_o | n6510_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6512_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n6514_o = n6512_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6515_o = n6511_o | n6514_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6516_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n6518_o = n6516_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6519_o = n6515_o | n6518_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6520_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n6522_o = n6520_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6523_o = n6519_o | n6522_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6524_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n6526_o = n6524_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6527_o = n6523_o | n6526_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6528_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n6530_o = n6528_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6531_o = n6527_o | n6530_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6532_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n6534_o = n6532_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6535_o = n6531_o | n6534_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6536_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n6538_o = n6536_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6539_o = n6535_o | n6538_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6540_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n6542_o = n6540_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6543_o = n6539_o | n6542_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6544_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n6546_o = n6544_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6547_o = n6543_o | n6546_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6548_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n6550_o = n6548_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6551_o = n6547_o | n6550_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6552_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n6554_o = n6552_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6555_o = n6551_o | n6554_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6556_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n6558_o = n6556_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6559_o = n6555_o | n6558_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6560_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n6562_o = n6560_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6563_o = n6559_o | n6562_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6564_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n6566_o = n6564_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6567_o = n6563_o | n6566_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6568_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n6570_o = n6568_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6571_o = n6567_o | n6570_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6572_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n6574_o = n6572_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6575_o = n6571_o | n6574_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6576_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n6578_o = n6576_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6579_o = n6575_o | n6578_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6580_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n6582_o = n6580_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6583_o = n6579_o | n6582_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6584_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n6586_o = n6584_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6587_o = n6583_o | n6586_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n6588_o = ~n6587_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n6589_o = ~n6588_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6601_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n6603_o = n6601_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6605_o = 1'b0 | n6603_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6607_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n6609_o = n6607_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6610_o = n6605_o | n6609_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6611_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n6613_o = n6611_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6614_o = n6610_o | n6613_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6615_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n6617_o = n6615_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6618_o = n6614_o | n6617_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6619_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n6621_o = n6619_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6622_o = n6618_o | n6621_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6623_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n6625_o = n6623_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6626_o = n6622_o | n6625_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6627_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n6629_o = n6627_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6630_o = n6626_o | n6629_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6631_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n6633_o = n6631_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6634_o = n6630_o | n6633_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6635_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n6637_o = n6635_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6638_o = n6634_o | n6637_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6639_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n6641_o = n6639_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6642_o = n6638_o | n6641_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6643_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n6645_o = n6643_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6646_o = n6642_o | n6645_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6647_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n6649_o = n6647_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6650_o = n6646_o | n6649_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6651_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n6653_o = n6651_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6654_o = n6650_o | n6653_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6655_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n6657_o = n6655_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6658_o = n6654_o | n6657_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6659_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n6661_o = n6659_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6662_o = n6658_o | n6661_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6663_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n6665_o = n6663_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6666_o = n6662_o | n6665_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6667_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n6669_o = n6667_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6670_o = n6666_o | n6669_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6671_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n6673_o = n6671_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6674_o = n6670_o | n6673_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6675_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n6677_o = n6675_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6678_o = n6674_o | n6677_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6679_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n6681_o = n6679_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6682_o = n6678_o | n6681_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6683_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n6685_o = n6683_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6686_o = n6682_o | n6685_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6687_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n6689_o = n6687_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6690_o = n6686_o | n6689_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6691_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n6693_o = n6691_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6694_o = n6690_o | n6693_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6695_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n6697_o = n6695_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6698_o = n6694_o | n6697_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6699_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n6701_o = n6699_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6702_o = n6698_o | n6701_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6703_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n6705_o = n6703_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6706_o = n6702_o | n6705_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6707_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n6709_o = n6707_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6710_o = n6706_o | n6709_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6711_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n6713_o = n6711_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6714_o = n6710_o | n6713_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6715_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n6717_o = n6715_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6718_o = n6714_o | n6717_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6719_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n6721_o = n6719_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6722_o = n6718_o | n6721_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6723_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n6725_o = n6723_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6726_o = n6722_o | n6725_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6727_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n6729_o = n6727_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6730_o = n6726_o | n6729_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n6731_o = ~n6730_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n6732_o = ~n6731_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6744_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n6746_o = n6744_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6748_o = 1'b0 | n6746_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6750_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n6752_o = n6750_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6753_o = n6748_o | n6752_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6754_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n6756_o = n6754_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6757_o = n6753_o | n6756_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6758_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n6760_o = n6758_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6761_o = n6757_o | n6760_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6762_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n6764_o = n6762_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6765_o = n6761_o | n6764_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6766_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n6768_o = n6766_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6769_o = n6765_o | n6768_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6770_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n6772_o = n6770_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6773_o = n6769_o | n6772_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6774_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n6776_o = n6774_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6777_o = n6773_o | n6776_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6778_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n6780_o = n6778_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6781_o = n6777_o | n6780_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6782_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n6784_o = n6782_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6785_o = n6781_o | n6784_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6786_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n6788_o = n6786_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6789_o = n6785_o | n6788_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6790_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n6792_o = n6790_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6793_o = n6789_o | n6792_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6794_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n6796_o = n6794_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6797_o = n6793_o | n6796_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6798_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n6800_o = n6798_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6801_o = n6797_o | n6800_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6802_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n6804_o = n6802_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6805_o = n6801_o | n6804_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6806_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n6808_o = n6806_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6809_o = n6805_o | n6808_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6810_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n6812_o = n6810_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6813_o = n6809_o | n6812_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6814_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n6816_o = n6814_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6817_o = n6813_o | n6816_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6818_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n6820_o = n6818_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6821_o = n6817_o | n6820_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6822_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n6824_o = n6822_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6825_o = n6821_o | n6824_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6826_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n6828_o = n6826_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6829_o = n6825_o | n6828_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6830_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n6832_o = n6830_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6833_o = n6829_o | n6832_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6834_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n6836_o = n6834_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6837_o = n6833_o | n6836_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6838_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n6840_o = n6838_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6841_o = n6837_o | n6840_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6842_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n6844_o = n6842_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6845_o = n6841_o | n6844_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6846_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n6848_o = n6846_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6849_o = n6845_o | n6848_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6850_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n6852_o = n6850_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6853_o = n6849_o | n6852_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6854_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n6856_o = n6854_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6857_o = n6853_o | n6856_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6858_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n6860_o = n6858_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6861_o = n6857_o | n6860_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6862_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n6864_o = n6862_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6865_o = n6861_o | n6864_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6866_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n6868_o = n6866_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6869_o = n6865_o | n6868_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6870_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n6872_o = n6870_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6873_o = n6869_o | n6872_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n6874_o = ~n6873_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n6875_o = ~n6874_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6887_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n6889_o = n6887_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6891_o = 1'b0 | n6889_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6893_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n6895_o = n6893_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6896_o = n6891_o | n6895_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6897_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n6899_o = n6897_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6900_o = n6896_o | n6899_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6901_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n6903_o = n6901_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6904_o = n6900_o | n6903_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6905_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n6907_o = n6905_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6908_o = n6904_o | n6907_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6909_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n6911_o = n6909_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6912_o = n6908_o | n6911_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6913_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n6915_o = n6913_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6916_o = n6912_o | n6915_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6917_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n6919_o = n6917_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6920_o = n6916_o | n6919_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6921_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n6923_o = n6921_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6924_o = n6920_o | n6923_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6925_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n6927_o = n6925_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6928_o = n6924_o | n6927_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6929_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n6931_o = n6929_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6932_o = n6928_o | n6931_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6933_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n6935_o = n6933_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6936_o = n6932_o | n6935_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6937_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n6939_o = n6937_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6940_o = n6936_o | n6939_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6941_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n6943_o = n6941_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6944_o = n6940_o | n6943_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6945_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n6947_o = n6945_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6948_o = n6944_o | n6947_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6949_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n6951_o = n6949_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6952_o = n6948_o | n6951_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6953_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n6955_o = n6953_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6956_o = n6952_o | n6955_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6957_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n6959_o = n6957_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6960_o = n6956_o | n6959_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6961_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n6963_o = n6961_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6964_o = n6960_o | n6963_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6965_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n6967_o = n6965_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6968_o = n6964_o | n6967_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6969_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n6971_o = n6969_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6972_o = n6968_o | n6971_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6973_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n6975_o = n6973_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6976_o = n6972_o | n6975_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6977_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n6979_o = n6977_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6980_o = n6976_o | n6979_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6981_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n6983_o = n6981_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n6984_o = n6980_o | n6983_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6985_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n6987_o = n6985_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6988_o = n6984_o | n6987_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6989_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n6991_o = n6989_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6992_o = n6988_o | n6991_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6993_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n6995_o = n6993_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n6996_o = n6992_o | n6995_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n6997_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n6999_o = n6997_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7000_o = n6996_o | n6999_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7001_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n7003_o = n7001_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7004_o = n7000_o | n7003_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7005_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n7007_o = n7005_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7008_o = n7004_o | n7007_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7009_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n7011_o = n7009_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7012_o = n7008_o | n7011_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7013_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n7015_o = n7013_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7016_o = n7012_o | n7015_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n7017_o = ~n7016_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n7018_o = ~n7017_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7030_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n7032_o = n7030_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7034_o = 1'b0 | n7032_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7036_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n7038_o = n7036_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7039_o = n7034_o | n7038_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7040_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n7042_o = n7040_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7043_o = n7039_o | n7042_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7044_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n7046_o = n7044_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7047_o = n7043_o | n7046_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7048_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n7050_o = n7048_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7051_o = n7047_o | n7050_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7052_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n7054_o = n7052_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7055_o = n7051_o | n7054_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7056_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n7058_o = n7056_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7059_o = n7055_o | n7058_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7060_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n7062_o = n7060_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7063_o = n7059_o | n7062_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7064_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n7066_o = n7064_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7067_o = n7063_o | n7066_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7068_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n7070_o = n7068_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7071_o = n7067_o | n7070_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7072_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n7074_o = n7072_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7075_o = n7071_o | n7074_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7076_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n7078_o = n7076_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7079_o = n7075_o | n7078_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7080_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n7082_o = n7080_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7083_o = n7079_o | n7082_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7084_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n7086_o = n7084_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7087_o = n7083_o | n7086_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7088_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n7090_o = n7088_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7091_o = n7087_o | n7090_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7092_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n7094_o = n7092_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7095_o = n7091_o | n7094_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7096_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n7098_o = n7096_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7099_o = n7095_o | n7098_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7100_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n7102_o = n7100_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7103_o = n7099_o | n7102_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7104_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n7106_o = n7104_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7107_o = n7103_o | n7106_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7108_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n7110_o = n7108_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7111_o = n7107_o | n7110_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7112_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n7114_o = n7112_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7115_o = n7111_o | n7114_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7116_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n7118_o = n7116_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7119_o = n7115_o | n7118_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7120_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n7122_o = n7120_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7123_o = n7119_o | n7122_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7124_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n7126_o = n7124_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7127_o = n7123_o | n7126_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7128_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n7130_o = n7128_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7131_o = n7127_o | n7130_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7132_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n7134_o = n7132_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7135_o = n7131_o | n7134_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7136_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n7138_o = n7136_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7139_o = n7135_o | n7138_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7140_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n7142_o = n7140_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7143_o = n7139_o | n7142_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7144_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n7146_o = n7144_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7147_o = n7143_o | n7146_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7148_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n7150_o = n7148_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7151_o = n7147_o | n7150_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7152_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n7154_o = n7152_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7155_o = n7151_o | n7154_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7156_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n7158_o = n7156_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7159_o = n7155_o | n7158_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n7160_o = ~n7159_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n7161_o = ~n7160_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7173_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n7175_o = n7173_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7177_o = 1'b0 | n7175_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7179_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n7181_o = n7179_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7182_o = n7177_o | n7181_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7183_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n7185_o = n7183_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7186_o = n7182_o | n7185_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7187_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n7189_o = n7187_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7190_o = n7186_o | n7189_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7191_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n7193_o = n7191_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7194_o = n7190_o | n7193_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7195_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n7197_o = n7195_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7198_o = n7194_o | n7197_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7199_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n7201_o = n7199_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7202_o = n7198_o | n7201_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7203_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n7205_o = n7203_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7206_o = n7202_o | n7205_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7207_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n7209_o = n7207_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7210_o = n7206_o | n7209_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7211_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n7213_o = n7211_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7214_o = n7210_o | n7213_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7215_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n7217_o = n7215_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7218_o = n7214_o | n7217_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7219_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n7221_o = n7219_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7222_o = n7218_o | n7221_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7223_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n7225_o = n7223_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7226_o = n7222_o | n7225_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7227_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n7229_o = n7227_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7230_o = n7226_o | n7229_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7231_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n7233_o = n7231_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7234_o = n7230_o | n7233_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7235_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n7237_o = n7235_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7238_o = n7234_o | n7237_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7239_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n7241_o = n7239_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7242_o = n7238_o | n7241_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7243_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n7245_o = n7243_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7246_o = n7242_o | n7245_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7247_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n7249_o = n7247_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7250_o = n7246_o | n7249_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7251_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n7253_o = n7251_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7254_o = n7250_o | n7253_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7255_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n7257_o = n7255_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7258_o = n7254_o | n7257_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7259_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n7261_o = n7259_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7262_o = n7258_o | n7261_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7263_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n7265_o = n7263_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7266_o = n7262_o | n7265_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7267_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n7269_o = n7267_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7270_o = n7266_o | n7269_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7271_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n7273_o = n7271_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7274_o = n7270_o | n7273_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7275_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n7277_o = n7275_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7278_o = n7274_o | n7277_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7279_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n7281_o = n7279_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7282_o = n7278_o | n7281_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7283_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n7285_o = n7283_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7286_o = n7282_o | n7285_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7287_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n7289_o = n7287_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7290_o = n7286_o | n7289_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7291_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n7293_o = n7291_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7294_o = n7290_o | n7293_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7295_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n7297_o = n7295_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7298_o = n7294_o | n7297_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7299_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n7301_o = n7299_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7302_o = n7298_o | n7301_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n7303_o = ~n7302_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n7304_o = ~n7303_o;
  assign n7305_o = {n7304_o, n7161_o, n7018_o, n6875_o};
  assign n7306_o = {n6732_o, n6589_o, n6446_o, n6303_o};
  assign n7307_o = {n6160_o, n6017_o};
  assign n7308_o = {n7305_o, n7306_o, n7307_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n7320_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n7322_o = n7320_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7324_o = 1'b0 | n7322_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7326_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n7328_o = n7326_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7329_o = n7324_o | n7328_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7330_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n7332_o = n7330_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7333_o = n7329_o | n7332_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7334_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n7336_o = n7334_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7337_o = n7333_o | n7336_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7338_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n7340_o = n7338_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7341_o = n7337_o | n7340_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7342_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n7344_o = n7342_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7345_o = n7341_o | n7344_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7346_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n7348_o = n7346_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7349_o = n7345_o | n7348_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7350_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n7352_o = n7350_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7353_o = n7349_o | n7352_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7354_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n7356_o = n7354_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7357_o = n7353_o | n7356_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7358_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n7360_o = n7358_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7361_o = n7357_o | n7360_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7362_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n7364_o = n7362_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7365_o = n7361_o | n7364_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7366_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n7368_o = n7366_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7369_o = n7365_o | n7368_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7370_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n7372_o = n7370_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7373_o = n7369_o | n7372_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7374_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n7376_o = n7374_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7377_o = n7373_o | n7376_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7378_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n7380_o = n7378_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7381_o = n7377_o | n7380_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7382_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n7384_o = n7382_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7385_o = n7381_o | n7384_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7386_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n7388_o = n7386_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7389_o = n7385_o | n7388_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7390_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n7392_o = n7390_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7393_o = n7389_o | n7392_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7394_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n7396_o = n7394_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7397_o = n7393_o | n7396_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7398_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n7400_o = n7398_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7401_o = n7397_o | n7400_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7402_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n7404_o = n7402_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7405_o = n7401_o | n7404_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7406_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n7408_o = n7406_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7409_o = n7405_o | n7408_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7410_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n7412_o = n7410_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7413_o = n7409_o | n7412_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7414_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n7416_o = n7414_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7417_o = n7413_o | n7416_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7418_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n7420_o = n7418_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7421_o = n7417_o | n7420_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7422_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n7424_o = n7422_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7425_o = n7421_o | n7424_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7426_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n7428_o = n7426_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7429_o = n7425_o | n7428_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7430_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n7432_o = n7430_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7433_o = n7429_o | n7432_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7434_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n7436_o = n7434_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7437_o = n7433_o | n7436_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7438_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n7440_o = n7438_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7441_o = n7437_o | n7440_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7442_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n7444_o = n7442_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7445_o = n7441_o | n7444_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7446_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n7448_o = n7446_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7449_o = n7445_o | n7448_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n7450_o = ~n7449_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n7451_o = ~n7450_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7463_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n7465_o = n7463_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7467_o = 1'b0 | n7465_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7469_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n7471_o = n7469_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7472_o = n7467_o | n7471_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7473_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n7475_o = n7473_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7476_o = n7472_o | n7475_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7477_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n7479_o = n7477_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7480_o = n7476_o | n7479_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7481_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n7483_o = n7481_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7484_o = n7480_o | n7483_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7485_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n7487_o = n7485_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7488_o = n7484_o | n7487_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7489_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n7491_o = n7489_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7492_o = n7488_o | n7491_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7493_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n7495_o = n7493_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7496_o = n7492_o | n7495_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7497_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n7499_o = n7497_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7500_o = n7496_o | n7499_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7501_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n7503_o = n7501_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7504_o = n7500_o | n7503_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7505_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n7507_o = n7505_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7508_o = n7504_o | n7507_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7509_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n7511_o = n7509_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7512_o = n7508_o | n7511_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7513_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n7515_o = n7513_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7516_o = n7512_o | n7515_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7517_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n7519_o = n7517_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7520_o = n7516_o | n7519_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7521_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n7523_o = n7521_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7524_o = n7520_o | n7523_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7525_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n7527_o = n7525_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7528_o = n7524_o | n7527_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7529_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n7531_o = n7529_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7532_o = n7528_o | n7531_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7533_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n7535_o = n7533_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7536_o = n7532_o | n7535_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7537_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n7539_o = n7537_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7540_o = n7536_o | n7539_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7541_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n7543_o = n7541_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7544_o = n7540_o | n7543_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7545_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n7547_o = n7545_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7548_o = n7544_o | n7547_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7549_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n7551_o = n7549_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7552_o = n7548_o | n7551_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7553_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n7555_o = n7553_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7556_o = n7552_o | n7555_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7557_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n7559_o = n7557_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7560_o = n7556_o | n7559_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7561_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n7563_o = n7561_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7564_o = n7560_o | n7563_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7565_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n7567_o = n7565_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7568_o = n7564_o | n7567_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7569_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n7571_o = n7569_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7572_o = n7568_o | n7571_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7573_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n7575_o = n7573_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7576_o = n7572_o | n7575_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7577_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n7579_o = n7577_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7580_o = n7576_o | n7579_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7581_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n7583_o = n7581_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7584_o = n7580_o | n7583_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7585_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n7587_o = n7585_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7588_o = n7584_o | n7587_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7589_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n7591_o = n7589_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7592_o = n7588_o | n7591_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n7593_o = ~n7592_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n7594_o = ~n7593_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7606_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n7608_o = n7606_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7610_o = 1'b0 | n7608_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7612_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n7614_o = n7612_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7615_o = n7610_o | n7614_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7616_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n7618_o = n7616_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7619_o = n7615_o | n7618_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7620_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n7622_o = n7620_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7623_o = n7619_o | n7622_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7624_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n7626_o = n7624_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7627_o = n7623_o | n7626_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7628_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n7630_o = n7628_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7631_o = n7627_o | n7630_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7632_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n7634_o = n7632_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7635_o = n7631_o | n7634_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7636_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n7638_o = n7636_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7639_o = n7635_o | n7638_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7640_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n7642_o = n7640_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7643_o = n7639_o | n7642_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7644_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n7646_o = n7644_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7647_o = n7643_o | n7646_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7648_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n7650_o = n7648_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7651_o = n7647_o | n7650_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7652_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n7654_o = n7652_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7655_o = n7651_o | n7654_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7656_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n7658_o = n7656_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7659_o = n7655_o | n7658_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7660_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n7662_o = n7660_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7663_o = n7659_o | n7662_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7664_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n7666_o = n7664_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7667_o = n7663_o | n7666_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7668_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n7670_o = n7668_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7671_o = n7667_o | n7670_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7672_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n7674_o = n7672_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7675_o = n7671_o | n7674_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7676_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n7678_o = n7676_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7679_o = n7675_o | n7678_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7680_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n7682_o = n7680_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7683_o = n7679_o | n7682_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7684_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n7686_o = n7684_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7687_o = n7683_o | n7686_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7688_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n7690_o = n7688_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7691_o = n7687_o | n7690_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7692_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n7694_o = n7692_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7695_o = n7691_o | n7694_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7696_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n7698_o = n7696_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7699_o = n7695_o | n7698_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7700_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n7702_o = n7700_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7703_o = n7699_o | n7702_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7704_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n7706_o = n7704_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7707_o = n7703_o | n7706_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7708_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n7710_o = n7708_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7711_o = n7707_o | n7710_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7712_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n7714_o = n7712_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7715_o = n7711_o | n7714_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7716_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n7718_o = n7716_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7719_o = n7715_o | n7718_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7720_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n7722_o = n7720_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7723_o = n7719_o | n7722_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7724_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n7726_o = n7724_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7727_o = n7723_o | n7726_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7728_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n7730_o = n7728_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7731_o = n7727_o | n7730_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7732_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n7734_o = n7732_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7735_o = n7731_o | n7734_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n7736_o = ~n7735_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n7737_o = ~n7736_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7749_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n7751_o = n7749_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7753_o = 1'b0 | n7751_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7755_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n7757_o = n7755_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7758_o = n7753_o | n7757_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7759_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n7761_o = n7759_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7762_o = n7758_o | n7761_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7763_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n7765_o = n7763_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7766_o = n7762_o | n7765_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7767_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n7769_o = n7767_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7770_o = n7766_o | n7769_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7771_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n7773_o = n7771_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7774_o = n7770_o | n7773_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7775_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n7777_o = n7775_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7778_o = n7774_o | n7777_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7779_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n7781_o = n7779_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7782_o = n7778_o | n7781_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7783_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n7785_o = n7783_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7786_o = n7782_o | n7785_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7787_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n7789_o = n7787_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7790_o = n7786_o | n7789_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7791_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n7793_o = n7791_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7794_o = n7790_o | n7793_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7795_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n7797_o = n7795_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7798_o = n7794_o | n7797_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7799_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n7801_o = n7799_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7802_o = n7798_o | n7801_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7803_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n7805_o = n7803_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7806_o = n7802_o | n7805_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7807_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n7809_o = n7807_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7810_o = n7806_o | n7809_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7811_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n7813_o = n7811_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7814_o = n7810_o | n7813_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7815_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n7817_o = n7815_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7818_o = n7814_o | n7817_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7819_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n7821_o = n7819_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7822_o = n7818_o | n7821_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7823_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n7825_o = n7823_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7826_o = n7822_o | n7825_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7827_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n7829_o = n7827_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7830_o = n7826_o | n7829_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7831_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n7833_o = n7831_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7834_o = n7830_o | n7833_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7835_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n7837_o = n7835_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7838_o = n7834_o | n7837_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7839_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n7841_o = n7839_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7842_o = n7838_o | n7841_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7843_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n7845_o = n7843_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7846_o = n7842_o | n7845_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7847_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n7849_o = n7847_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7850_o = n7846_o | n7849_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7851_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n7853_o = n7851_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7854_o = n7850_o | n7853_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7855_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n7857_o = n7855_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7858_o = n7854_o | n7857_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7859_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n7861_o = n7859_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7862_o = n7858_o | n7861_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7863_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n7865_o = n7863_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7866_o = n7862_o | n7865_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7867_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n7869_o = n7867_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7870_o = n7866_o | n7869_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7871_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n7873_o = n7871_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7874_o = n7870_o | n7873_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7875_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n7877_o = n7875_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7878_o = n7874_o | n7877_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n7879_o = ~n7878_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n7880_o = ~n7879_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7892_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n7894_o = n7892_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7896_o = 1'b0 | n7894_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7898_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n7900_o = n7898_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7901_o = n7896_o | n7900_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7902_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n7904_o = n7902_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7905_o = n7901_o | n7904_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7906_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n7908_o = n7906_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7909_o = n7905_o | n7908_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7910_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n7912_o = n7910_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7913_o = n7909_o | n7912_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7914_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n7916_o = n7914_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7917_o = n7913_o | n7916_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7918_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n7920_o = n7918_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7921_o = n7917_o | n7920_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7922_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n7924_o = n7922_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7925_o = n7921_o | n7924_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7926_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n7928_o = n7926_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7929_o = n7925_o | n7928_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7930_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n7932_o = n7930_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7933_o = n7929_o | n7932_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7934_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n7936_o = n7934_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7937_o = n7933_o | n7936_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7938_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n7940_o = n7938_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7941_o = n7937_o | n7940_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7942_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n7944_o = n7942_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7945_o = n7941_o | n7944_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7946_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n7948_o = n7946_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7949_o = n7945_o | n7948_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7950_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n7952_o = n7950_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7953_o = n7949_o | n7952_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7954_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n7956_o = n7954_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7957_o = n7953_o | n7956_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7958_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n7960_o = n7958_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7961_o = n7957_o | n7960_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7962_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n7964_o = n7962_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7965_o = n7961_o | n7964_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7966_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n7968_o = n7966_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7969_o = n7965_o | n7968_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7970_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n7972_o = n7970_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7973_o = n7969_o | n7972_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7974_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n7976_o = n7974_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7977_o = n7973_o | n7976_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7978_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n7980_o = n7978_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7981_o = n7977_o | n7980_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7982_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n7984_o = n7982_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7985_o = n7981_o | n7984_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7986_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n7988_o = n7986_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7989_o = n7985_o | n7988_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7990_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n7992_o = n7990_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n7993_o = n7989_o | n7992_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7994_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n7996_o = n7994_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n7997_o = n7993_o | n7996_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n7998_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n8000_o = n7998_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8001_o = n7997_o | n8000_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8002_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n8004_o = n8002_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8005_o = n8001_o | n8004_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8006_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n8008_o = n8006_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8009_o = n8005_o | n8008_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8010_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n8012_o = n8010_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8013_o = n8009_o | n8012_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8014_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n8016_o = n8014_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8017_o = n8013_o | n8016_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8018_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n8020_o = n8018_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8021_o = n8017_o | n8020_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n8022_o = ~n8021_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n8023_o = ~n8022_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8035_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n8037_o = n8035_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8039_o = 1'b0 | n8037_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8041_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n8043_o = n8041_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8044_o = n8039_o | n8043_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8045_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n8047_o = n8045_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8048_o = n8044_o | n8047_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8049_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n8051_o = n8049_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8052_o = n8048_o | n8051_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8053_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n8055_o = n8053_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8056_o = n8052_o | n8055_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8057_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n8059_o = n8057_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8060_o = n8056_o | n8059_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8061_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n8063_o = n8061_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8064_o = n8060_o | n8063_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8065_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n8067_o = n8065_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8068_o = n8064_o | n8067_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8069_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n8071_o = n8069_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8072_o = n8068_o | n8071_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8073_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n8075_o = n8073_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8076_o = n8072_o | n8075_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8077_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n8079_o = n8077_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8080_o = n8076_o | n8079_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8081_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n8083_o = n8081_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8084_o = n8080_o | n8083_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8085_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n8087_o = n8085_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8088_o = n8084_o | n8087_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8089_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n8091_o = n8089_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8092_o = n8088_o | n8091_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8093_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n8095_o = n8093_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8096_o = n8092_o | n8095_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8097_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n8099_o = n8097_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8100_o = n8096_o | n8099_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8101_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n8103_o = n8101_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8104_o = n8100_o | n8103_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8105_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n8107_o = n8105_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8108_o = n8104_o | n8107_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8109_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n8111_o = n8109_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8112_o = n8108_o | n8111_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8113_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n8115_o = n8113_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8116_o = n8112_o | n8115_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8117_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n8119_o = n8117_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8120_o = n8116_o | n8119_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8121_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n8123_o = n8121_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8124_o = n8120_o | n8123_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8125_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n8127_o = n8125_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8128_o = n8124_o | n8127_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8129_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n8131_o = n8129_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8132_o = n8128_o | n8131_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8133_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n8135_o = n8133_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8136_o = n8132_o | n8135_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8137_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n8139_o = n8137_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8140_o = n8136_o | n8139_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8141_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n8143_o = n8141_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8144_o = n8140_o | n8143_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8145_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n8147_o = n8145_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8148_o = n8144_o | n8147_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8149_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n8151_o = n8149_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8152_o = n8148_o | n8151_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8153_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n8155_o = n8153_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8156_o = n8152_o | n8155_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8157_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n8159_o = n8157_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8160_o = n8156_o | n8159_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8161_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n8163_o = n8161_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8164_o = n8160_o | n8163_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n8165_o = ~n8164_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n8166_o = ~n8165_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8178_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n8180_o = n8178_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8182_o = 1'b0 | n8180_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8184_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n8186_o = n8184_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8187_o = n8182_o | n8186_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8188_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n8190_o = n8188_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8191_o = n8187_o | n8190_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8192_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n8194_o = n8192_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8195_o = n8191_o | n8194_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8196_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n8198_o = n8196_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8199_o = n8195_o | n8198_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8200_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n8202_o = n8200_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8203_o = n8199_o | n8202_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8204_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n8206_o = n8204_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8207_o = n8203_o | n8206_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8208_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n8210_o = n8208_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8211_o = n8207_o | n8210_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8212_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n8214_o = n8212_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8215_o = n8211_o | n8214_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8216_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n8218_o = n8216_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8219_o = n8215_o | n8218_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8220_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n8222_o = n8220_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8223_o = n8219_o | n8222_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8224_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n8226_o = n8224_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8227_o = n8223_o | n8226_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8228_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n8230_o = n8228_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8231_o = n8227_o | n8230_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8232_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n8234_o = n8232_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8235_o = n8231_o | n8234_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8236_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n8238_o = n8236_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8239_o = n8235_o | n8238_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8240_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n8242_o = n8240_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8243_o = n8239_o | n8242_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8244_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n8246_o = n8244_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8247_o = n8243_o | n8246_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8248_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n8250_o = n8248_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8251_o = n8247_o | n8250_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8252_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n8254_o = n8252_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8255_o = n8251_o | n8254_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8256_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n8258_o = n8256_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8259_o = n8255_o | n8258_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8260_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n8262_o = n8260_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8263_o = n8259_o | n8262_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8264_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n8266_o = n8264_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8267_o = n8263_o | n8266_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8268_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n8270_o = n8268_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8271_o = n8267_o | n8270_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8272_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n8274_o = n8272_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8275_o = n8271_o | n8274_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8276_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n8278_o = n8276_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8279_o = n8275_o | n8278_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8280_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n8282_o = n8280_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8283_o = n8279_o | n8282_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8284_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n8286_o = n8284_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8287_o = n8283_o | n8286_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8288_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n8290_o = n8288_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8291_o = n8287_o | n8290_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8292_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n8294_o = n8292_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8295_o = n8291_o | n8294_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8296_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n8298_o = n8296_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8299_o = n8295_o | n8298_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8300_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n8302_o = n8300_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8303_o = n8299_o | n8302_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8304_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n8306_o = n8304_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8307_o = n8303_o | n8306_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n8308_o = ~n8307_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n8309_o = ~n8308_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8321_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n8323_o = n8321_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8325_o = 1'b0 | n8323_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8327_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n8329_o = n8327_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8330_o = n8325_o | n8329_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8331_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n8333_o = n8331_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8334_o = n8330_o | n8333_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8335_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n8337_o = n8335_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8338_o = n8334_o | n8337_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8339_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n8341_o = n8339_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8342_o = n8338_o | n8341_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8343_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n8345_o = n8343_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8346_o = n8342_o | n8345_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8347_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n8349_o = n8347_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8350_o = n8346_o | n8349_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8351_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n8353_o = n8351_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8354_o = n8350_o | n8353_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8355_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n8357_o = n8355_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8358_o = n8354_o | n8357_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8359_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n8361_o = n8359_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8362_o = n8358_o | n8361_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8363_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n8365_o = n8363_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8366_o = n8362_o | n8365_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8367_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n8369_o = n8367_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8370_o = n8366_o | n8369_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8371_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n8373_o = n8371_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8374_o = n8370_o | n8373_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8375_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n8377_o = n8375_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8378_o = n8374_o | n8377_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8379_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n8381_o = n8379_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8382_o = n8378_o | n8381_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8383_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n8385_o = n8383_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8386_o = n8382_o | n8385_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8387_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n8389_o = n8387_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8390_o = n8386_o | n8389_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8391_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n8393_o = n8391_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8394_o = n8390_o | n8393_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8395_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n8397_o = n8395_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8398_o = n8394_o | n8397_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8399_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n8401_o = n8399_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8402_o = n8398_o | n8401_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8403_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n8405_o = n8403_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8406_o = n8402_o | n8405_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8407_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n8409_o = n8407_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8410_o = n8406_o | n8409_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8411_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n8413_o = n8411_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8414_o = n8410_o | n8413_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8415_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n8417_o = n8415_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8418_o = n8414_o | n8417_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8419_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n8421_o = n8419_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8422_o = n8418_o | n8421_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8423_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n8425_o = n8423_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8426_o = n8422_o | n8425_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8427_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n8429_o = n8427_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8430_o = n8426_o | n8429_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8431_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n8433_o = n8431_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8434_o = n8430_o | n8433_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8435_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n8437_o = n8435_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8438_o = n8434_o | n8437_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8439_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n8441_o = n8439_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8442_o = n8438_o | n8441_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8443_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n8445_o = n8443_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8446_o = n8442_o | n8445_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8447_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n8449_o = n8447_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8450_o = n8446_o | n8449_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n8451_o = ~n8450_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n8452_o = ~n8451_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8464_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n8466_o = n8464_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8468_o = 1'b0 | n8466_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8470_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n8472_o = n8470_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8473_o = n8468_o | n8472_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8474_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n8476_o = n8474_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8477_o = n8473_o | n8476_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8478_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n8480_o = n8478_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8481_o = n8477_o | n8480_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8482_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n8484_o = n8482_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8485_o = n8481_o | n8484_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8486_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n8488_o = n8486_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8489_o = n8485_o | n8488_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8490_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n8492_o = n8490_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8493_o = n8489_o | n8492_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8494_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n8496_o = n8494_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8497_o = n8493_o | n8496_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8498_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n8500_o = n8498_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8501_o = n8497_o | n8500_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8502_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n8504_o = n8502_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8505_o = n8501_o | n8504_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8506_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n8508_o = n8506_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8509_o = n8505_o | n8508_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8510_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n8512_o = n8510_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8513_o = n8509_o | n8512_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8514_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n8516_o = n8514_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8517_o = n8513_o | n8516_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8518_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n8520_o = n8518_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8521_o = n8517_o | n8520_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8522_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n8524_o = n8522_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8525_o = n8521_o | n8524_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8526_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n8528_o = n8526_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8529_o = n8525_o | n8528_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8530_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n8532_o = n8530_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8533_o = n8529_o | n8532_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8534_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n8536_o = n8534_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8537_o = n8533_o | n8536_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8538_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n8540_o = n8538_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8541_o = n8537_o | n8540_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8542_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n8544_o = n8542_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8545_o = n8541_o | n8544_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8546_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n8548_o = n8546_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8549_o = n8545_o | n8548_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8550_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n8552_o = n8550_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8553_o = n8549_o | n8552_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8554_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n8556_o = n8554_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8557_o = n8553_o | n8556_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8558_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n8560_o = n8558_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8561_o = n8557_o | n8560_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8562_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n8564_o = n8562_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8565_o = n8561_o | n8564_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8566_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n8568_o = n8566_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8569_o = n8565_o | n8568_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8570_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n8572_o = n8570_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8573_o = n8569_o | n8572_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8574_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n8576_o = n8574_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8577_o = n8573_o | n8576_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8578_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n8580_o = n8578_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8581_o = n8577_o | n8580_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8582_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n8584_o = n8582_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8585_o = n8581_o | n8584_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8586_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n8588_o = n8586_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8589_o = n8585_o | n8588_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8590_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n8592_o = n8590_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8593_o = n8589_o | n8592_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n8594_o = ~n8593_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n8595_o = ~n8594_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8607_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n8609_o = n8607_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8611_o = 1'b0 | n8609_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8613_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n8615_o = n8613_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8616_o = n8611_o | n8615_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8617_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n8619_o = n8617_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8620_o = n8616_o | n8619_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8621_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n8623_o = n8621_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8624_o = n8620_o | n8623_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8625_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n8627_o = n8625_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8628_o = n8624_o | n8627_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8629_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n8631_o = n8629_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8632_o = n8628_o | n8631_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8633_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n8635_o = n8633_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8636_o = n8632_o | n8635_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8637_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n8639_o = n8637_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8640_o = n8636_o | n8639_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8641_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n8643_o = n8641_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8644_o = n8640_o | n8643_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8645_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n8647_o = n8645_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8648_o = n8644_o | n8647_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8649_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n8651_o = n8649_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8652_o = n8648_o | n8651_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8653_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n8655_o = n8653_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8656_o = n8652_o | n8655_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8657_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n8659_o = n8657_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8660_o = n8656_o | n8659_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8661_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n8663_o = n8661_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8664_o = n8660_o | n8663_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8665_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n8667_o = n8665_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8668_o = n8664_o | n8667_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8669_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n8671_o = n8669_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8672_o = n8668_o | n8671_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8673_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n8675_o = n8673_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8676_o = n8672_o | n8675_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8677_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n8679_o = n8677_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8680_o = n8676_o | n8679_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8681_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n8683_o = n8681_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8684_o = n8680_o | n8683_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8685_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n8687_o = n8685_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8688_o = n8684_o | n8687_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8689_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n8691_o = n8689_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8692_o = n8688_o | n8691_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8693_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n8695_o = n8693_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8696_o = n8692_o | n8695_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8697_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n8699_o = n8697_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8700_o = n8696_o | n8699_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8701_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n8703_o = n8701_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8704_o = n8700_o | n8703_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8705_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n8707_o = n8705_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8708_o = n8704_o | n8707_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8709_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n8711_o = n8709_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8712_o = n8708_o | n8711_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8713_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n8715_o = n8713_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8716_o = n8712_o | n8715_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8717_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n8719_o = n8717_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8720_o = n8716_o | n8719_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8721_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n8723_o = n8721_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8724_o = n8720_o | n8723_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8725_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n8727_o = n8725_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8728_o = n8724_o | n8727_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8729_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n8731_o = n8729_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8732_o = n8728_o | n8731_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8733_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n8735_o = n8733_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8736_o = n8732_o | n8735_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n8737_o = ~n8736_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n8738_o = ~n8737_o;
  assign n8739_o = {n8738_o, n8595_o, n8452_o, n8309_o};
  assign n8740_o = {n8166_o, n8023_o, n7880_o, n7737_o};
  assign n8741_o = {n7594_o, n7451_o};
  assign n8742_o = {n8739_o, n8740_o, n8741_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n8754_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n8756_o = n8754_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8758_o = 1'b0 | n8756_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8760_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n8762_o = n8760_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8763_o = n8758_o | n8762_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8764_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n8766_o = n8764_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8767_o = n8763_o | n8766_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8768_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n8770_o = n8768_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8771_o = n8767_o | n8770_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8772_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n8774_o = n8772_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8775_o = n8771_o | n8774_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8776_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n8778_o = n8776_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8779_o = n8775_o | n8778_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8780_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n8782_o = n8780_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8783_o = n8779_o | n8782_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8784_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n8786_o = n8784_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8787_o = n8783_o | n8786_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8788_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n8790_o = n8788_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8791_o = n8787_o | n8790_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8792_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n8794_o = n8792_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8795_o = n8791_o | n8794_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8796_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n8798_o = n8796_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8799_o = n8795_o | n8798_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8800_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n8802_o = n8800_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8803_o = n8799_o | n8802_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8804_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n8806_o = n8804_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8807_o = n8803_o | n8806_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8808_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n8810_o = n8808_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8811_o = n8807_o | n8810_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8812_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n8814_o = n8812_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8815_o = n8811_o | n8814_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8816_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n8818_o = n8816_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8819_o = n8815_o | n8818_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8820_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n8822_o = n8820_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8823_o = n8819_o | n8822_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8824_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n8826_o = n8824_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8827_o = n8823_o | n8826_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8828_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n8830_o = n8828_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8831_o = n8827_o | n8830_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8832_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n8834_o = n8832_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8835_o = n8831_o | n8834_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8836_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n8838_o = n8836_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8839_o = n8835_o | n8838_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8840_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n8842_o = n8840_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8843_o = n8839_o | n8842_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8844_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n8846_o = n8844_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8847_o = n8843_o | n8846_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8848_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n8850_o = n8848_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8851_o = n8847_o | n8850_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8852_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n8854_o = n8852_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8855_o = n8851_o | n8854_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8856_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n8858_o = n8856_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8859_o = n8855_o | n8858_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8860_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n8862_o = n8860_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8863_o = n8859_o | n8862_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8864_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n8866_o = n8864_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8867_o = n8863_o | n8866_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8868_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n8870_o = n8868_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8871_o = n8867_o | n8870_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8872_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n8874_o = n8872_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8875_o = n8871_o | n8874_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8876_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n8878_o = n8876_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8879_o = n8875_o | n8878_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8880_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n8882_o = n8880_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8883_o = n8879_o | n8882_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n8884_o = ~n8883_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n8885_o = ~n8884_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8897_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n8899_o = n8897_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8901_o = 1'b0 | n8899_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8903_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n8905_o = n8903_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8906_o = n8901_o | n8905_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8907_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n8909_o = n8907_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8910_o = n8906_o | n8909_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8911_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n8913_o = n8911_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8914_o = n8910_o | n8913_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8915_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n8917_o = n8915_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8918_o = n8914_o | n8917_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8919_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n8921_o = n8919_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8922_o = n8918_o | n8921_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8923_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n8925_o = n8923_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8926_o = n8922_o | n8925_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8927_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n8929_o = n8927_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8930_o = n8926_o | n8929_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8931_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n8933_o = n8931_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8934_o = n8930_o | n8933_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8935_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n8937_o = n8935_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8938_o = n8934_o | n8937_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8939_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n8941_o = n8939_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8942_o = n8938_o | n8941_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8943_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n8945_o = n8943_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8946_o = n8942_o | n8945_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8947_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n8949_o = n8947_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8950_o = n8946_o | n8949_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8951_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n8953_o = n8951_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8954_o = n8950_o | n8953_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8955_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n8957_o = n8955_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8958_o = n8954_o | n8957_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8959_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n8961_o = n8959_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8962_o = n8958_o | n8961_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8963_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n8965_o = n8963_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8966_o = n8962_o | n8965_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8967_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n8969_o = n8967_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8970_o = n8966_o | n8969_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8971_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n8973_o = n8971_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8974_o = n8970_o | n8973_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8975_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n8977_o = n8975_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8978_o = n8974_o | n8977_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8979_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n8981_o = n8979_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8982_o = n8978_o | n8981_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8983_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n8985_o = n8983_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8986_o = n8982_o | n8985_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8987_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n8989_o = n8987_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8990_o = n8986_o | n8989_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8991_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n8993_o = n8991_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n8994_o = n8990_o | n8993_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8995_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n8997_o = n8995_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n8998_o = n8994_o | n8997_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n8999_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n9001_o = n8999_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9002_o = n8998_o | n9001_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9003_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n9005_o = n9003_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9006_o = n9002_o | n9005_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9007_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n9009_o = n9007_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9010_o = n9006_o | n9009_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9011_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n9013_o = n9011_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9014_o = n9010_o | n9013_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9015_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n9017_o = n9015_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9018_o = n9014_o | n9017_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9019_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n9021_o = n9019_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9022_o = n9018_o | n9021_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9023_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n9025_o = n9023_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9026_o = n9022_o | n9025_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n9027_o = ~n9026_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n9028_o = ~n9027_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9040_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n9042_o = n9040_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9044_o = 1'b0 | n9042_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9046_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n9048_o = n9046_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9049_o = n9044_o | n9048_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9050_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n9052_o = n9050_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9053_o = n9049_o | n9052_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9054_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n9056_o = n9054_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9057_o = n9053_o | n9056_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9058_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n9060_o = n9058_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9061_o = n9057_o | n9060_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9062_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n9064_o = n9062_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9065_o = n9061_o | n9064_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9066_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n9068_o = n9066_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9069_o = n9065_o | n9068_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9070_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n9072_o = n9070_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9073_o = n9069_o | n9072_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9074_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n9076_o = n9074_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9077_o = n9073_o | n9076_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9078_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n9080_o = n9078_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9081_o = n9077_o | n9080_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9082_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n9084_o = n9082_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9085_o = n9081_o | n9084_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9086_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n9088_o = n9086_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9089_o = n9085_o | n9088_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9090_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n9092_o = n9090_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9093_o = n9089_o | n9092_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9094_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n9096_o = n9094_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9097_o = n9093_o | n9096_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9098_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n9100_o = n9098_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9101_o = n9097_o | n9100_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9102_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n9104_o = n9102_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9105_o = n9101_o | n9104_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9106_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n9108_o = n9106_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9109_o = n9105_o | n9108_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9110_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n9112_o = n9110_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9113_o = n9109_o | n9112_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9114_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n9116_o = n9114_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9117_o = n9113_o | n9116_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9118_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n9120_o = n9118_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9121_o = n9117_o | n9120_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9122_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n9124_o = n9122_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9125_o = n9121_o | n9124_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9126_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n9128_o = n9126_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9129_o = n9125_o | n9128_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9130_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n9132_o = n9130_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9133_o = n9129_o | n9132_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9134_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n9136_o = n9134_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9137_o = n9133_o | n9136_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9138_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n9140_o = n9138_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9141_o = n9137_o | n9140_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9142_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n9144_o = n9142_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9145_o = n9141_o | n9144_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9146_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n9148_o = n9146_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9149_o = n9145_o | n9148_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9150_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n9152_o = n9150_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9153_o = n9149_o | n9152_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9154_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n9156_o = n9154_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9157_o = n9153_o | n9156_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9158_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n9160_o = n9158_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9161_o = n9157_o | n9160_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9162_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n9164_o = n9162_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9165_o = n9161_o | n9164_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9166_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n9168_o = n9166_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9169_o = n9165_o | n9168_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n9170_o = ~n9169_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n9171_o = ~n9170_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9183_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n9185_o = n9183_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9187_o = 1'b0 | n9185_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9189_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n9191_o = n9189_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9192_o = n9187_o | n9191_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9193_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n9195_o = n9193_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9196_o = n9192_o | n9195_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9197_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n9199_o = n9197_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9200_o = n9196_o | n9199_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9201_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n9203_o = n9201_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9204_o = n9200_o | n9203_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9205_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n9207_o = n9205_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9208_o = n9204_o | n9207_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9209_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n9211_o = n9209_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9212_o = n9208_o | n9211_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9213_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n9215_o = n9213_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9216_o = n9212_o | n9215_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9217_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n9219_o = n9217_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9220_o = n9216_o | n9219_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9221_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n9223_o = n9221_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9224_o = n9220_o | n9223_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9225_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n9227_o = n9225_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9228_o = n9224_o | n9227_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9229_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n9231_o = n9229_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9232_o = n9228_o | n9231_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9233_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n9235_o = n9233_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9236_o = n9232_o | n9235_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9237_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n9239_o = n9237_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9240_o = n9236_o | n9239_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9241_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n9243_o = n9241_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9244_o = n9240_o | n9243_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9245_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n9247_o = n9245_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9248_o = n9244_o | n9247_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9249_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n9251_o = n9249_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9252_o = n9248_o | n9251_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9253_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n9255_o = n9253_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9256_o = n9252_o | n9255_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9257_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n9259_o = n9257_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9260_o = n9256_o | n9259_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9261_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n9263_o = n9261_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9264_o = n9260_o | n9263_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9265_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n9267_o = n9265_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9268_o = n9264_o | n9267_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9269_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n9271_o = n9269_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9272_o = n9268_o | n9271_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9273_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n9275_o = n9273_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9276_o = n9272_o | n9275_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9277_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n9279_o = n9277_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9280_o = n9276_o | n9279_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9281_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n9283_o = n9281_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9284_o = n9280_o | n9283_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9285_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n9287_o = n9285_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9288_o = n9284_o | n9287_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9289_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n9291_o = n9289_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9292_o = n9288_o | n9291_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9293_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n9295_o = n9293_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9296_o = n9292_o | n9295_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9297_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n9299_o = n9297_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9300_o = n9296_o | n9299_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9301_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n9303_o = n9301_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9304_o = n9300_o | n9303_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9305_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n9307_o = n9305_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9308_o = n9304_o | n9307_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9309_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n9311_o = n9309_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9312_o = n9308_o | n9311_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n9313_o = ~n9312_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n9314_o = ~n9313_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9326_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n9328_o = n9326_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9330_o = 1'b0 | n9328_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9332_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n9334_o = n9332_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9335_o = n9330_o | n9334_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9336_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n9338_o = n9336_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9339_o = n9335_o | n9338_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9340_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n9342_o = n9340_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9343_o = n9339_o | n9342_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9344_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n9346_o = n9344_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9347_o = n9343_o | n9346_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9348_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n9350_o = n9348_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9351_o = n9347_o | n9350_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9352_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n9354_o = n9352_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9355_o = n9351_o | n9354_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9356_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n9358_o = n9356_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9359_o = n9355_o | n9358_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9360_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n9362_o = n9360_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9363_o = n9359_o | n9362_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9364_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n9366_o = n9364_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9367_o = n9363_o | n9366_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9368_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n9370_o = n9368_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9371_o = n9367_o | n9370_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9372_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n9374_o = n9372_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9375_o = n9371_o | n9374_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9376_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n9378_o = n9376_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9379_o = n9375_o | n9378_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9380_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n9382_o = n9380_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9383_o = n9379_o | n9382_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9384_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n9386_o = n9384_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9387_o = n9383_o | n9386_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9388_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n9390_o = n9388_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9391_o = n9387_o | n9390_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9392_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n9394_o = n9392_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9395_o = n9391_o | n9394_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9396_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n9398_o = n9396_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9399_o = n9395_o | n9398_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9400_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n9402_o = n9400_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9403_o = n9399_o | n9402_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9404_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n9406_o = n9404_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9407_o = n9403_o | n9406_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9408_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n9410_o = n9408_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9411_o = n9407_o | n9410_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9412_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n9414_o = n9412_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9415_o = n9411_o | n9414_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9416_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n9418_o = n9416_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9419_o = n9415_o | n9418_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9420_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n9422_o = n9420_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9423_o = n9419_o | n9422_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9424_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n9426_o = n9424_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9427_o = n9423_o | n9426_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9428_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n9430_o = n9428_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9431_o = n9427_o | n9430_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9432_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n9434_o = n9432_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9435_o = n9431_o | n9434_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9436_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n9438_o = n9436_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9439_o = n9435_o | n9438_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9440_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n9442_o = n9440_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9443_o = n9439_o | n9442_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9444_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n9446_o = n9444_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9447_o = n9443_o | n9446_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9448_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n9450_o = n9448_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9451_o = n9447_o | n9450_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9452_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n9454_o = n9452_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9455_o = n9451_o | n9454_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n9456_o = ~n9455_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n9457_o = ~n9456_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9469_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n9471_o = n9469_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9473_o = 1'b0 | n9471_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9475_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n9477_o = n9475_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9478_o = n9473_o | n9477_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9479_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n9481_o = n9479_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9482_o = n9478_o | n9481_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9483_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n9485_o = n9483_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9486_o = n9482_o | n9485_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9487_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n9489_o = n9487_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9490_o = n9486_o | n9489_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9491_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n9493_o = n9491_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9494_o = n9490_o | n9493_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9495_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n9497_o = n9495_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9498_o = n9494_o | n9497_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9499_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n9501_o = n9499_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9502_o = n9498_o | n9501_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9503_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n9505_o = n9503_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9506_o = n9502_o | n9505_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9507_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n9509_o = n9507_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9510_o = n9506_o | n9509_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9511_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n9513_o = n9511_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9514_o = n9510_o | n9513_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9515_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n9517_o = n9515_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9518_o = n9514_o | n9517_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9519_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n9521_o = n9519_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9522_o = n9518_o | n9521_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9523_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n9525_o = n9523_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9526_o = n9522_o | n9525_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9527_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n9529_o = n9527_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9530_o = n9526_o | n9529_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9531_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n9533_o = n9531_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9534_o = n9530_o | n9533_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9535_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n9537_o = n9535_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9538_o = n9534_o | n9537_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9539_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n9541_o = n9539_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9542_o = n9538_o | n9541_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9543_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n9545_o = n9543_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9546_o = n9542_o | n9545_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9547_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n9549_o = n9547_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9550_o = n9546_o | n9549_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9551_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n9553_o = n9551_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9554_o = n9550_o | n9553_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9555_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n9557_o = n9555_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9558_o = n9554_o | n9557_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9559_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n9561_o = n9559_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9562_o = n9558_o | n9561_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9563_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n9565_o = n9563_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9566_o = n9562_o | n9565_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9567_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n9569_o = n9567_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9570_o = n9566_o | n9569_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9571_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n9573_o = n9571_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9574_o = n9570_o | n9573_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9575_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n9577_o = n9575_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9578_o = n9574_o | n9577_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9579_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n9581_o = n9579_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9582_o = n9578_o | n9581_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9583_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n9585_o = n9583_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9586_o = n9582_o | n9585_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9587_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n9589_o = n9587_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9590_o = n9586_o | n9589_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9591_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n9593_o = n9591_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9594_o = n9590_o | n9593_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9595_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n9597_o = n9595_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9598_o = n9594_o | n9597_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n9599_o = ~n9598_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n9600_o = ~n9599_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9612_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n9614_o = n9612_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9616_o = 1'b0 | n9614_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9618_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n9620_o = n9618_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9621_o = n9616_o | n9620_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9622_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n9624_o = n9622_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9625_o = n9621_o | n9624_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9626_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n9628_o = n9626_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9629_o = n9625_o | n9628_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9630_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n9632_o = n9630_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9633_o = n9629_o | n9632_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9634_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n9636_o = n9634_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9637_o = n9633_o | n9636_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9638_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n9640_o = n9638_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9641_o = n9637_o | n9640_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9642_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n9644_o = n9642_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9645_o = n9641_o | n9644_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9646_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n9648_o = n9646_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9649_o = n9645_o | n9648_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9650_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n9652_o = n9650_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9653_o = n9649_o | n9652_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9654_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n9656_o = n9654_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9657_o = n9653_o | n9656_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9658_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n9660_o = n9658_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9661_o = n9657_o | n9660_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9662_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n9664_o = n9662_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9665_o = n9661_o | n9664_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9666_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n9668_o = n9666_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9669_o = n9665_o | n9668_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9670_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n9672_o = n9670_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9673_o = n9669_o | n9672_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9674_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n9676_o = n9674_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9677_o = n9673_o | n9676_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9678_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n9680_o = n9678_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9681_o = n9677_o | n9680_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9682_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n9684_o = n9682_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9685_o = n9681_o | n9684_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9686_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n9688_o = n9686_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9689_o = n9685_o | n9688_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9690_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n9692_o = n9690_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9693_o = n9689_o | n9692_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9694_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n9696_o = n9694_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9697_o = n9693_o | n9696_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9698_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n9700_o = n9698_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9701_o = n9697_o | n9700_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9702_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n9704_o = n9702_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9705_o = n9701_o | n9704_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9706_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n9708_o = n9706_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9709_o = n9705_o | n9708_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9710_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n9712_o = n9710_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9713_o = n9709_o | n9712_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9714_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n9716_o = n9714_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9717_o = n9713_o | n9716_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9718_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n9720_o = n9718_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9721_o = n9717_o | n9720_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9722_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n9724_o = n9722_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9725_o = n9721_o | n9724_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9726_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n9728_o = n9726_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9729_o = n9725_o | n9728_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9730_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n9732_o = n9730_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9733_o = n9729_o | n9732_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9734_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n9736_o = n9734_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9737_o = n9733_o | n9736_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9738_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n9740_o = n9738_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9741_o = n9737_o | n9740_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n9742_o = ~n9741_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n9743_o = ~n9742_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9755_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n9757_o = n9755_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9759_o = 1'b0 | n9757_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9761_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n9763_o = n9761_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9764_o = n9759_o | n9763_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9765_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n9767_o = n9765_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9768_o = n9764_o | n9767_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9769_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n9771_o = n9769_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9772_o = n9768_o | n9771_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9773_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n9775_o = n9773_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9776_o = n9772_o | n9775_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9777_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n9779_o = n9777_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9780_o = n9776_o | n9779_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9781_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n9783_o = n9781_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9784_o = n9780_o | n9783_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9785_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n9787_o = n9785_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9788_o = n9784_o | n9787_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9789_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n9791_o = n9789_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9792_o = n9788_o | n9791_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9793_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n9795_o = n9793_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9796_o = n9792_o | n9795_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9797_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n9799_o = n9797_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9800_o = n9796_o | n9799_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9801_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n9803_o = n9801_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9804_o = n9800_o | n9803_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9805_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n9807_o = n9805_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9808_o = n9804_o | n9807_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9809_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n9811_o = n9809_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9812_o = n9808_o | n9811_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9813_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n9815_o = n9813_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9816_o = n9812_o | n9815_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9817_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n9819_o = n9817_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9820_o = n9816_o | n9819_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9821_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n9823_o = n9821_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9824_o = n9820_o | n9823_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9825_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n9827_o = n9825_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9828_o = n9824_o | n9827_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9829_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n9831_o = n9829_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9832_o = n9828_o | n9831_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9833_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n9835_o = n9833_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9836_o = n9832_o | n9835_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9837_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n9839_o = n9837_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9840_o = n9836_o | n9839_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9841_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n9843_o = n9841_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9844_o = n9840_o | n9843_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9845_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n9847_o = n9845_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9848_o = n9844_o | n9847_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9849_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n9851_o = n9849_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9852_o = n9848_o | n9851_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9853_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n9855_o = n9853_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9856_o = n9852_o | n9855_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9857_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n9859_o = n9857_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9860_o = n9856_o | n9859_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9861_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n9863_o = n9861_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9864_o = n9860_o | n9863_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9865_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n9867_o = n9865_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9868_o = n9864_o | n9867_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9869_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n9871_o = n9869_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9872_o = n9868_o | n9871_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9873_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n9875_o = n9873_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9876_o = n9872_o | n9875_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9877_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n9879_o = n9877_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9880_o = n9876_o | n9879_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9881_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n9883_o = n9881_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9884_o = n9880_o | n9883_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n9885_o = ~n9884_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n9886_o = ~n9885_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9898_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n9900_o = n9898_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9902_o = 1'b0 | n9900_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9904_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n9906_o = n9904_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9907_o = n9902_o | n9906_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9908_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n9910_o = n9908_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9911_o = n9907_o | n9910_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9912_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n9914_o = n9912_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9915_o = n9911_o | n9914_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9916_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n9918_o = n9916_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9919_o = n9915_o | n9918_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9920_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n9922_o = n9920_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9923_o = n9919_o | n9922_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9924_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n9926_o = n9924_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9927_o = n9923_o | n9926_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9928_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n9930_o = n9928_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9931_o = n9927_o | n9930_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9932_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n9934_o = n9932_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9935_o = n9931_o | n9934_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9936_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n9938_o = n9936_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9939_o = n9935_o | n9938_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9940_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n9942_o = n9940_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9943_o = n9939_o | n9942_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9944_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n9946_o = n9944_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9947_o = n9943_o | n9946_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9948_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n9950_o = n9948_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9951_o = n9947_o | n9950_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9952_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n9954_o = n9952_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9955_o = n9951_o | n9954_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9956_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n9958_o = n9956_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9959_o = n9955_o | n9958_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9960_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n9962_o = n9960_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n9963_o = n9959_o | n9962_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9964_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n9966_o = n9964_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9967_o = n9963_o | n9966_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9968_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n9970_o = n9968_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9971_o = n9967_o | n9970_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9972_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n9974_o = n9972_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9975_o = n9971_o | n9974_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9976_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n9978_o = n9976_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9979_o = n9975_o | n9978_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9980_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n9982_o = n9980_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9983_o = n9979_o | n9982_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9984_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n9986_o = n9984_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9987_o = n9983_o | n9986_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9988_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n9990_o = n9988_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9991_o = n9987_o | n9990_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9992_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n9994_o = n9992_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9995_o = n9991_o | n9994_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n9996_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n9998_o = n9996_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n9999_o = n9995_o | n9998_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10000_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n10002_o = n10000_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10003_o = n9999_o | n10002_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10004_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n10006_o = n10004_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10007_o = n10003_o | n10006_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10008_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n10010_o = n10008_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10011_o = n10007_o | n10010_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10012_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n10014_o = n10012_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10015_o = n10011_o | n10014_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10016_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n10018_o = n10016_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10019_o = n10015_o | n10018_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10020_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n10022_o = n10020_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10023_o = n10019_o | n10022_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10024_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n10026_o = n10024_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10027_o = n10023_o | n10026_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n10028_o = ~n10027_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n10029_o = ~n10028_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10041_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n10043_o = n10041_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10045_o = 1'b0 | n10043_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10047_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n10049_o = n10047_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10050_o = n10045_o | n10049_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10051_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n10053_o = n10051_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10054_o = n10050_o | n10053_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10055_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n10057_o = n10055_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10058_o = n10054_o | n10057_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10059_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n10061_o = n10059_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10062_o = n10058_o | n10061_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10063_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n10065_o = n10063_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10066_o = n10062_o | n10065_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10067_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n10069_o = n10067_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10070_o = n10066_o | n10069_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10071_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n10073_o = n10071_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10074_o = n10070_o | n10073_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10075_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n10077_o = n10075_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10078_o = n10074_o | n10077_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10079_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n10081_o = n10079_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10082_o = n10078_o | n10081_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10083_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n10085_o = n10083_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10086_o = n10082_o | n10085_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10087_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n10089_o = n10087_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10090_o = n10086_o | n10089_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10091_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n10093_o = n10091_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10094_o = n10090_o | n10093_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10095_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n10097_o = n10095_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10098_o = n10094_o | n10097_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10099_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n10101_o = n10099_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10102_o = n10098_o | n10101_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10103_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n10105_o = n10103_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10106_o = n10102_o | n10105_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10107_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n10109_o = n10107_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10110_o = n10106_o | n10109_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10111_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n10113_o = n10111_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10114_o = n10110_o | n10113_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10115_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n10117_o = n10115_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10118_o = n10114_o | n10117_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10119_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n10121_o = n10119_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10122_o = n10118_o | n10121_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10123_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n10125_o = n10123_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10126_o = n10122_o | n10125_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10127_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n10129_o = n10127_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10130_o = n10126_o | n10129_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10131_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n10133_o = n10131_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10134_o = n10130_o | n10133_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10135_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n10137_o = n10135_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10138_o = n10134_o | n10137_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10139_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n10141_o = n10139_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10142_o = n10138_o | n10141_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10143_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n10145_o = n10143_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10146_o = n10142_o | n10145_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10147_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n10149_o = n10147_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10150_o = n10146_o | n10149_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10151_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n10153_o = n10151_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10154_o = n10150_o | n10153_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10155_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n10157_o = n10155_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10158_o = n10154_o | n10157_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10159_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n10161_o = n10159_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10162_o = n10158_o | n10161_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10163_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n10165_o = n10163_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10166_o = n10162_o | n10165_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10167_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n10169_o = n10167_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10170_o = n10166_o | n10169_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n10171_o = ~n10170_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n10172_o = ~n10171_o;
  assign n10173_o = {n10172_o, n10029_o, n9886_o, n9743_o};
  assign n10174_o = {n9600_o, n9457_o, n9314_o, n9171_o};
  assign n10175_o = {n9028_o, n8885_o};
  assign n10176_o = {n10173_o, n10174_o, n10175_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n10188_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n10190_o = n10188_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10192_o = 1'b0 | n10190_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10194_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n10196_o = n10194_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10197_o = n10192_o | n10196_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10198_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n10200_o = n10198_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10201_o = n10197_o | n10200_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10202_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n10204_o = n10202_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10205_o = n10201_o | n10204_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10206_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n10208_o = n10206_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10209_o = n10205_o | n10208_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10210_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n10212_o = n10210_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10213_o = n10209_o | n10212_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10214_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n10216_o = n10214_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10217_o = n10213_o | n10216_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10218_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n10220_o = n10218_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10221_o = n10217_o | n10220_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10222_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n10224_o = n10222_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10225_o = n10221_o | n10224_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10226_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n10228_o = n10226_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10229_o = n10225_o | n10228_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10230_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n10232_o = n10230_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10233_o = n10229_o | n10232_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10234_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n10236_o = n10234_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10237_o = n10233_o | n10236_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10238_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n10240_o = n10238_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10241_o = n10237_o | n10240_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10242_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n10244_o = n10242_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10245_o = n10241_o | n10244_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10246_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n10248_o = n10246_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10249_o = n10245_o | n10248_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10250_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n10252_o = n10250_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10253_o = n10249_o | n10252_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10254_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n10256_o = n10254_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10257_o = n10253_o | n10256_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10258_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n10260_o = n10258_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10261_o = n10257_o | n10260_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10262_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n10264_o = n10262_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10265_o = n10261_o | n10264_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10266_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n10268_o = n10266_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10269_o = n10265_o | n10268_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10270_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n10272_o = n10270_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10273_o = n10269_o | n10272_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10274_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n10276_o = n10274_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10277_o = n10273_o | n10276_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10278_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n10280_o = n10278_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10281_o = n10277_o | n10280_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10282_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n10284_o = n10282_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10285_o = n10281_o | n10284_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10286_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n10288_o = n10286_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10289_o = n10285_o | n10288_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10290_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n10292_o = n10290_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10293_o = n10289_o | n10292_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10294_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n10296_o = n10294_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10297_o = n10293_o | n10296_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10298_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n10300_o = n10298_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10301_o = n10297_o | n10300_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10302_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n10304_o = n10302_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10305_o = n10301_o | n10304_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10306_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n10308_o = n10306_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10309_o = n10305_o | n10308_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10310_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n10312_o = n10310_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10313_o = n10309_o | n10312_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10314_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n10316_o = n10314_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10317_o = n10313_o | n10316_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n10318_o = ~n10317_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n10319_o = ~n10318_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10331_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n10333_o = n10331_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10335_o = 1'b0 | n10333_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10337_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n10339_o = n10337_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10340_o = n10335_o | n10339_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10341_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n10343_o = n10341_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10344_o = n10340_o | n10343_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10345_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n10347_o = n10345_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10348_o = n10344_o | n10347_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10349_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n10351_o = n10349_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10352_o = n10348_o | n10351_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10353_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n10355_o = n10353_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10356_o = n10352_o | n10355_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10357_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n10359_o = n10357_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10360_o = n10356_o | n10359_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10361_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n10363_o = n10361_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10364_o = n10360_o | n10363_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10365_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n10367_o = n10365_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10368_o = n10364_o | n10367_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10369_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n10371_o = n10369_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10372_o = n10368_o | n10371_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10373_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n10375_o = n10373_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10376_o = n10372_o | n10375_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10377_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n10379_o = n10377_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10380_o = n10376_o | n10379_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10381_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n10383_o = n10381_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10384_o = n10380_o | n10383_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10385_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n10387_o = n10385_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10388_o = n10384_o | n10387_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10389_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n10391_o = n10389_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10392_o = n10388_o | n10391_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10393_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n10395_o = n10393_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10396_o = n10392_o | n10395_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10397_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n10399_o = n10397_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10400_o = n10396_o | n10399_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10401_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n10403_o = n10401_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10404_o = n10400_o | n10403_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10405_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n10407_o = n10405_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10408_o = n10404_o | n10407_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10409_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n10411_o = n10409_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10412_o = n10408_o | n10411_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10413_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n10415_o = n10413_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10416_o = n10412_o | n10415_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10417_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n10419_o = n10417_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10420_o = n10416_o | n10419_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10421_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n10423_o = n10421_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10424_o = n10420_o | n10423_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10425_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n10427_o = n10425_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10428_o = n10424_o | n10427_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10429_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n10431_o = n10429_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10432_o = n10428_o | n10431_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10433_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n10435_o = n10433_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10436_o = n10432_o | n10435_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10437_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n10439_o = n10437_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10440_o = n10436_o | n10439_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10441_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n10443_o = n10441_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10444_o = n10440_o | n10443_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10445_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n10447_o = n10445_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10448_o = n10444_o | n10447_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10449_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n10451_o = n10449_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10452_o = n10448_o | n10451_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10453_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n10455_o = n10453_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10456_o = n10452_o | n10455_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10457_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n10459_o = n10457_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10460_o = n10456_o | n10459_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n10461_o = ~n10460_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n10462_o = ~n10461_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10474_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n10476_o = n10474_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10478_o = 1'b0 | n10476_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10480_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n10482_o = n10480_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10483_o = n10478_o | n10482_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10484_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n10486_o = n10484_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10487_o = n10483_o | n10486_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10488_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n10490_o = n10488_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10491_o = n10487_o | n10490_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10492_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n10494_o = n10492_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10495_o = n10491_o | n10494_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10496_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n10498_o = n10496_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10499_o = n10495_o | n10498_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10500_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n10502_o = n10500_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10503_o = n10499_o | n10502_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10504_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n10506_o = n10504_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10507_o = n10503_o | n10506_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10508_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n10510_o = n10508_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10511_o = n10507_o | n10510_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10512_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n10514_o = n10512_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10515_o = n10511_o | n10514_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10516_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n10518_o = n10516_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10519_o = n10515_o | n10518_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10520_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n10522_o = n10520_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10523_o = n10519_o | n10522_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10524_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n10526_o = n10524_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10527_o = n10523_o | n10526_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10528_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n10530_o = n10528_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10531_o = n10527_o | n10530_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10532_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n10534_o = n10532_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10535_o = n10531_o | n10534_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10536_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n10538_o = n10536_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10539_o = n10535_o | n10538_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10540_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n10542_o = n10540_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10543_o = n10539_o | n10542_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10544_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n10546_o = n10544_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10547_o = n10543_o | n10546_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10548_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n10550_o = n10548_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10551_o = n10547_o | n10550_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10552_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n10554_o = n10552_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10555_o = n10551_o | n10554_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10556_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n10558_o = n10556_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10559_o = n10555_o | n10558_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10560_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n10562_o = n10560_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10563_o = n10559_o | n10562_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10564_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n10566_o = n10564_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10567_o = n10563_o | n10566_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10568_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n10570_o = n10568_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10571_o = n10567_o | n10570_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10572_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n10574_o = n10572_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10575_o = n10571_o | n10574_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10576_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n10578_o = n10576_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10579_o = n10575_o | n10578_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10580_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n10582_o = n10580_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10583_o = n10579_o | n10582_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10584_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n10586_o = n10584_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10587_o = n10583_o | n10586_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10588_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n10590_o = n10588_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10591_o = n10587_o | n10590_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10592_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n10594_o = n10592_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10595_o = n10591_o | n10594_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10596_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n10598_o = n10596_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10599_o = n10595_o | n10598_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10600_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n10602_o = n10600_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10603_o = n10599_o | n10602_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n10604_o = ~n10603_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n10605_o = ~n10604_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10617_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n10619_o = n10617_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10621_o = 1'b0 | n10619_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10623_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n10625_o = n10623_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10626_o = n10621_o | n10625_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10627_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n10629_o = n10627_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10630_o = n10626_o | n10629_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10631_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n10633_o = n10631_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10634_o = n10630_o | n10633_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10635_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n10637_o = n10635_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10638_o = n10634_o | n10637_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10639_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n10641_o = n10639_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10642_o = n10638_o | n10641_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10643_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n10645_o = n10643_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10646_o = n10642_o | n10645_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10647_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n10649_o = n10647_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10650_o = n10646_o | n10649_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10651_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n10653_o = n10651_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10654_o = n10650_o | n10653_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10655_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n10657_o = n10655_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10658_o = n10654_o | n10657_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10659_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n10661_o = n10659_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10662_o = n10658_o | n10661_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10663_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n10665_o = n10663_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10666_o = n10662_o | n10665_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10667_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n10669_o = n10667_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10670_o = n10666_o | n10669_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10671_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n10673_o = n10671_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10674_o = n10670_o | n10673_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10675_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n10677_o = n10675_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10678_o = n10674_o | n10677_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10679_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n10681_o = n10679_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10682_o = n10678_o | n10681_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10683_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n10685_o = n10683_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10686_o = n10682_o | n10685_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10687_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n10689_o = n10687_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10690_o = n10686_o | n10689_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10691_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n10693_o = n10691_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10694_o = n10690_o | n10693_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10695_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n10697_o = n10695_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10698_o = n10694_o | n10697_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10699_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n10701_o = n10699_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10702_o = n10698_o | n10701_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10703_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n10705_o = n10703_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10706_o = n10702_o | n10705_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10707_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n10709_o = n10707_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10710_o = n10706_o | n10709_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10711_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n10713_o = n10711_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10714_o = n10710_o | n10713_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10715_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n10717_o = n10715_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10718_o = n10714_o | n10717_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10719_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n10721_o = n10719_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10722_o = n10718_o | n10721_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10723_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n10725_o = n10723_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10726_o = n10722_o | n10725_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10727_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n10729_o = n10727_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10730_o = n10726_o | n10729_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10731_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n10733_o = n10731_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10734_o = n10730_o | n10733_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10735_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n10737_o = n10735_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10738_o = n10734_o | n10737_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10739_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n10741_o = n10739_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10742_o = n10738_o | n10741_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10743_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n10745_o = n10743_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10746_o = n10742_o | n10745_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n10747_o = ~n10746_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n10748_o = ~n10747_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10760_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n10762_o = n10760_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10764_o = 1'b0 | n10762_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10766_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n10768_o = n10766_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10769_o = n10764_o | n10768_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10770_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n10772_o = n10770_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10773_o = n10769_o | n10772_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10774_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n10776_o = n10774_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10777_o = n10773_o | n10776_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10778_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n10780_o = n10778_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10781_o = n10777_o | n10780_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10782_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n10784_o = n10782_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10785_o = n10781_o | n10784_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10786_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n10788_o = n10786_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10789_o = n10785_o | n10788_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10790_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n10792_o = n10790_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10793_o = n10789_o | n10792_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10794_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n10796_o = n10794_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10797_o = n10793_o | n10796_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10798_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n10800_o = n10798_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10801_o = n10797_o | n10800_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10802_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n10804_o = n10802_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10805_o = n10801_o | n10804_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10806_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n10808_o = n10806_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10809_o = n10805_o | n10808_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10810_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n10812_o = n10810_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10813_o = n10809_o | n10812_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10814_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n10816_o = n10814_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10817_o = n10813_o | n10816_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10818_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n10820_o = n10818_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10821_o = n10817_o | n10820_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10822_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n10824_o = n10822_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10825_o = n10821_o | n10824_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10826_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n10828_o = n10826_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10829_o = n10825_o | n10828_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10830_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n10832_o = n10830_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10833_o = n10829_o | n10832_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10834_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n10836_o = n10834_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10837_o = n10833_o | n10836_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10838_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n10840_o = n10838_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10841_o = n10837_o | n10840_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10842_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n10844_o = n10842_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10845_o = n10841_o | n10844_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10846_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n10848_o = n10846_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10849_o = n10845_o | n10848_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10850_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n10852_o = n10850_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10853_o = n10849_o | n10852_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10854_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n10856_o = n10854_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10857_o = n10853_o | n10856_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10858_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n10860_o = n10858_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10861_o = n10857_o | n10860_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10862_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n10864_o = n10862_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10865_o = n10861_o | n10864_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10866_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n10868_o = n10866_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10869_o = n10865_o | n10868_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10870_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n10872_o = n10870_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10873_o = n10869_o | n10872_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10874_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n10876_o = n10874_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10877_o = n10873_o | n10876_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10878_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n10880_o = n10878_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10881_o = n10877_o | n10880_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10882_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n10884_o = n10882_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10885_o = n10881_o | n10884_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10886_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n10888_o = n10886_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10889_o = n10885_o | n10888_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n10890_o = ~n10889_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n10891_o = ~n10890_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10903_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n10905_o = n10903_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10907_o = 1'b0 | n10905_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10909_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n10911_o = n10909_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10912_o = n10907_o | n10911_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10913_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n10915_o = n10913_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10916_o = n10912_o | n10915_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10917_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n10919_o = n10917_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10920_o = n10916_o | n10919_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10921_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n10923_o = n10921_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10924_o = n10920_o | n10923_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10925_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n10927_o = n10925_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10928_o = n10924_o | n10927_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10929_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n10931_o = n10929_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10932_o = n10928_o | n10931_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10933_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n10935_o = n10933_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10936_o = n10932_o | n10935_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10937_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n10939_o = n10937_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10940_o = n10936_o | n10939_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10941_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n10943_o = n10941_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10944_o = n10940_o | n10943_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10945_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n10947_o = n10945_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10948_o = n10944_o | n10947_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10949_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n10951_o = n10949_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10952_o = n10948_o | n10951_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10953_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n10955_o = n10953_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10956_o = n10952_o | n10955_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10957_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n10959_o = n10957_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10960_o = n10956_o | n10959_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10961_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n10963_o = n10961_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10964_o = n10960_o | n10963_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10965_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n10967_o = n10965_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10968_o = n10964_o | n10967_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10969_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n10971_o = n10969_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n10972_o = n10968_o | n10971_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10973_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n10975_o = n10973_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10976_o = n10972_o | n10975_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10977_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n10979_o = n10977_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10980_o = n10976_o | n10979_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10981_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n10983_o = n10981_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10984_o = n10980_o | n10983_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10985_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n10987_o = n10985_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10988_o = n10984_o | n10987_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10989_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n10991_o = n10989_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10992_o = n10988_o | n10991_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10993_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n10995_o = n10993_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n10996_o = n10992_o | n10995_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n10997_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n10999_o = n10997_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11000_o = n10996_o | n10999_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11001_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n11003_o = n11001_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11004_o = n11000_o | n11003_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11005_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n11007_o = n11005_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11008_o = n11004_o | n11007_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11009_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n11011_o = n11009_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11012_o = n11008_o | n11011_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11013_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n11015_o = n11013_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11016_o = n11012_o | n11015_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11017_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n11019_o = n11017_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11020_o = n11016_o | n11019_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11021_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n11023_o = n11021_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11024_o = n11020_o | n11023_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11025_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n11027_o = n11025_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11028_o = n11024_o | n11027_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11029_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n11031_o = n11029_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11032_o = n11028_o | n11031_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n11033_o = ~n11032_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n11034_o = ~n11033_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11046_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n11048_o = n11046_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11050_o = 1'b0 | n11048_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11052_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n11054_o = n11052_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11055_o = n11050_o | n11054_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11056_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n11058_o = n11056_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11059_o = n11055_o | n11058_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11060_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n11062_o = n11060_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11063_o = n11059_o | n11062_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11064_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n11066_o = n11064_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11067_o = n11063_o | n11066_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11068_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n11070_o = n11068_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11071_o = n11067_o | n11070_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11072_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n11074_o = n11072_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11075_o = n11071_o | n11074_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11076_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n11078_o = n11076_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11079_o = n11075_o | n11078_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11080_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n11082_o = n11080_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11083_o = n11079_o | n11082_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11084_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n11086_o = n11084_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11087_o = n11083_o | n11086_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11088_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n11090_o = n11088_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11091_o = n11087_o | n11090_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11092_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n11094_o = n11092_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11095_o = n11091_o | n11094_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11096_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n11098_o = n11096_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11099_o = n11095_o | n11098_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11100_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n11102_o = n11100_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11103_o = n11099_o | n11102_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11104_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n11106_o = n11104_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11107_o = n11103_o | n11106_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11108_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n11110_o = n11108_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11111_o = n11107_o | n11110_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11112_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n11114_o = n11112_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11115_o = n11111_o | n11114_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11116_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n11118_o = n11116_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11119_o = n11115_o | n11118_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11120_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n11122_o = n11120_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11123_o = n11119_o | n11122_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11124_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n11126_o = n11124_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11127_o = n11123_o | n11126_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11128_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n11130_o = n11128_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11131_o = n11127_o | n11130_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11132_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n11134_o = n11132_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11135_o = n11131_o | n11134_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11136_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n11138_o = n11136_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11139_o = n11135_o | n11138_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11140_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n11142_o = n11140_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11143_o = n11139_o | n11142_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11144_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n11146_o = n11144_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11147_o = n11143_o | n11146_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11148_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n11150_o = n11148_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11151_o = n11147_o | n11150_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11152_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n11154_o = n11152_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11155_o = n11151_o | n11154_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11156_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n11158_o = n11156_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11159_o = n11155_o | n11158_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11160_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n11162_o = n11160_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11163_o = n11159_o | n11162_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11164_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n11166_o = n11164_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11167_o = n11163_o | n11166_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11168_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n11170_o = n11168_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11171_o = n11167_o | n11170_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11172_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n11174_o = n11172_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11175_o = n11171_o | n11174_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n11176_o = ~n11175_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n11177_o = ~n11176_o;
  assign n11181_o = {1'b0, 1'b0, 1'b0, n11177_o};
  assign n11182_o = {n11034_o, n10891_o, n10748_o, n10605_o};
  assign n11183_o = {n10462_o, n10319_o};
  assign n11184_o = {n11181_o, n11182_o, n11183_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n11196_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n11198_o = n11196_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11200_o = 1'b0 | n11198_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11202_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n11204_o = n11202_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11205_o = n11200_o | n11204_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11206_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n11208_o = n11206_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11209_o = n11205_o | n11208_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11210_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n11212_o = n11210_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11213_o = n11209_o | n11212_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11214_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n11216_o = n11214_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11217_o = n11213_o | n11216_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11218_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n11220_o = n11218_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11221_o = n11217_o | n11220_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11222_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n11224_o = n11222_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11225_o = n11221_o | n11224_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11226_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n11228_o = n11226_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11229_o = n11225_o | n11228_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11230_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n11232_o = n11230_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11233_o = n11229_o | n11232_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11234_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n11236_o = n11234_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11237_o = n11233_o | n11236_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11238_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n11240_o = n11238_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11241_o = n11237_o | n11240_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11242_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n11244_o = n11242_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11245_o = n11241_o | n11244_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11246_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n11248_o = n11246_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11249_o = n11245_o | n11248_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11250_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n11252_o = n11250_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11253_o = n11249_o | n11252_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11254_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n11256_o = n11254_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11257_o = n11253_o | n11256_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11258_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n11260_o = n11258_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11261_o = n11257_o | n11260_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11262_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n11264_o = n11262_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11265_o = n11261_o | n11264_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11266_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n11268_o = n11266_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11269_o = n11265_o | n11268_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11270_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n11272_o = n11270_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11273_o = n11269_o | n11272_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11274_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n11276_o = n11274_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11277_o = n11273_o | n11276_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11278_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n11280_o = n11278_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11281_o = n11277_o | n11280_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11282_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n11284_o = n11282_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11285_o = n11281_o | n11284_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11286_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n11288_o = n11286_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11289_o = n11285_o | n11288_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11290_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n11292_o = n11290_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11293_o = n11289_o | n11292_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11294_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n11296_o = n11294_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11297_o = n11293_o | n11296_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11298_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n11300_o = n11298_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11301_o = n11297_o | n11300_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11302_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n11304_o = n11302_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11305_o = n11301_o | n11304_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11306_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n11308_o = n11306_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11309_o = n11305_o | n11308_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11310_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n11312_o = n11310_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11313_o = n11309_o | n11312_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11314_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n11316_o = n11314_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11317_o = n11313_o | n11316_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11318_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n11320_o = n11318_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11321_o = n11317_o | n11320_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11322_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n11324_o = n11322_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11325_o = n11321_o | n11324_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n11326_o = ~n11325_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n11327_o = ~n11326_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11339_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n11341_o = n11339_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11343_o = 1'b0 | n11341_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11345_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n11347_o = n11345_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11348_o = n11343_o | n11347_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11349_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n11351_o = n11349_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11352_o = n11348_o | n11351_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11353_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n11355_o = n11353_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11356_o = n11352_o | n11355_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11357_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n11359_o = n11357_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11360_o = n11356_o | n11359_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11361_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n11363_o = n11361_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11364_o = n11360_o | n11363_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11365_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n11367_o = n11365_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11368_o = n11364_o | n11367_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11369_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n11371_o = n11369_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11372_o = n11368_o | n11371_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11373_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n11375_o = n11373_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11376_o = n11372_o | n11375_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11377_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n11379_o = n11377_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11380_o = n11376_o | n11379_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11381_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n11383_o = n11381_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11384_o = n11380_o | n11383_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11385_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n11387_o = n11385_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11388_o = n11384_o | n11387_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11389_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n11391_o = n11389_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11392_o = n11388_o | n11391_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11393_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n11395_o = n11393_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11396_o = n11392_o | n11395_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11397_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n11399_o = n11397_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11400_o = n11396_o | n11399_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11401_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n11403_o = n11401_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11404_o = n11400_o | n11403_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11405_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n11407_o = n11405_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11408_o = n11404_o | n11407_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11409_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n11411_o = n11409_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11412_o = n11408_o | n11411_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11413_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n11415_o = n11413_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11416_o = n11412_o | n11415_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11417_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n11419_o = n11417_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11420_o = n11416_o | n11419_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11421_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n11423_o = n11421_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11424_o = n11420_o | n11423_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11425_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n11427_o = n11425_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11428_o = n11424_o | n11427_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11429_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n11431_o = n11429_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11432_o = n11428_o | n11431_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11433_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n11435_o = n11433_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11436_o = n11432_o | n11435_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11437_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n11439_o = n11437_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11440_o = n11436_o | n11439_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11441_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n11443_o = n11441_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11444_o = n11440_o | n11443_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11445_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n11447_o = n11445_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11448_o = n11444_o | n11447_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11449_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n11451_o = n11449_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11452_o = n11448_o | n11451_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11453_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n11455_o = n11453_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11456_o = n11452_o | n11455_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11457_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n11459_o = n11457_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11460_o = n11456_o | n11459_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11461_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n11463_o = n11461_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11464_o = n11460_o | n11463_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11465_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n11467_o = n11465_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11468_o = n11464_o | n11467_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n11469_o = ~n11468_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n11470_o = ~n11469_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11482_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n11484_o = n11482_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11486_o = 1'b0 | n11484_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11488_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n11490_o = n11488_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11491_o = n11486_o | n11490_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11492_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n11494_o = n11492_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11495_o = n11491_o | n11494_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11496_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n11498_o = n11496_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11499_o = n11495_o | n11498_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11500_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n11502_o = n11500_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11503_o = n11499_o | n11502_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11504_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n11506_o = n11504_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11507_o = n11503_o | n11506_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11508_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n11510_o = n11508_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11511_o = n11507_o | n11510_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11512_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n11514_o = n11512_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11515_o = n11511_o | n11514_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11516_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n11518_o = n11516_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11519_o = n11515_o | n11518_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11520_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n11522_o = n11520_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11523_o = n11519_o | n11522_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11524_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n11526_o = n11524_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11527_o = n11523_o | n11526_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11528_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n11530_o = n11528_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11531_o = n11527_o | n11530_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11532_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n11534_o = n11532_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11535_o = n11531_o | n11534_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11536_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n11538_o = n11536_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11539_o = n11535_o | n11538_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11540_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n11542_o = n11540_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11543_o = n11539_o | n11542_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11544_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n11546_o = n11544_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11547_o = n11543_o | n11546_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11548_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n11550_o = n11548_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11551_o = n11547_o | n11550_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11552_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n11554_o = n11552_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11555_o = n11551_o | n11554_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11556_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n11558_o = n11556_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11559_o = n11555_o | n11558_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11560_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n11562_o = n11560_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11563_o = n11559_o | n11562_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11564_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n11566_o = n11564_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11567_o = n11563_o | n11566_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11568_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n11570_o = n11568_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11571_o = n11567_o | n11570_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11572_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n11574_o = n11572_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11575_o = n11571_o | n11574_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11576_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n11578_o = n11576_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11579_o = n11575_o | n11578_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11580_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n11582_o = n11580_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11583_o = n11579_o | n11582_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11584_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n11586_o = n11584_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11587_o = n11583_o | n11586_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11588_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n11590_o = n11588_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11591_o = n11587_o | n11590_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11592_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n11594_o = n11592_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11595_o = n11591_o | n11594_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11596_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n11598_o = n11596_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11599_o = n11595_o | n11598_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11600_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n11602_o = n11600_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11603_o = n11599_o | n11602_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11604_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n11606_o = n11604_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11607_o = n11603_o | n11606_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11608_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n11610_o = n11608_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11611_o = n11607_o | n11610_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n11612_o = ~n11611_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n11613_o = ~n11612_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11625_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n11627_o = n11625_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11629_o = 1'b0 | n11627_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11631_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n11633_o = n11631_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11634_o = n11629_o | n11633_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11635_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n11637_o = n11635_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11638_o = n11634_o | n11637_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11639_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n11641_o = n11639_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11642_o = n11638_o | n11641_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11643_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n11645_o = n11643_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11646_o = n11642_o | n11645_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11647_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n11649_o = n11647_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11650_o = n11646_o | n11649_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11651_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n11653_o = n11651_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11654_o = n11650_o | n11653_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11655_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n11657_o = n11655_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11658_o = n11654_o | n11657_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11659_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n11661_o = n11659_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11662_o = n11658_o | n11661_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11663_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n11665_o = n11663_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11666_o = n11662_o | n11665_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11667_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n11669_o = n11667_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11670_o = n11666_o | n11669_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11671_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n11673_o = n11671_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11674_o = n11670_o | n11673_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11675_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n11677_o = n11675_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11678_o = n11674_o | n11677_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11679_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n11681_o = n11679_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11682_o = n11678_o | n11681_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11683_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n11685_o = n11683_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11686_o = n11682_o | n11685_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11687_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n11689_o = n11687_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11690_o = n11686_o | n11689_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11691_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n11693_o = n11691_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11694_o = n11690_o | n11693_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11695_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n11697_o = n11695_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11698_o = n11694_o | n11697_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11699_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n11701_o = n11699_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11702_o = n11698_o | n11701_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11703_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n11705_o = n11703_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11706_o = n11702_o | n11705_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11707_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n11709_o = n11707_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11710_o = n11706_o | n11709_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11711_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n11713_o = n11711_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11714_o = n11710_o | n11713_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11715_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n11717_o = n11715_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11718_o = n11714_o | n11717_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11719_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n11721_o = n11719_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11722_o = n11718_o | n11721_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11723_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n11725_o = n11723_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11726_o = n11722_o | n11725_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11727_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n11729_o = n11727_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11730_o = n11726_o | n11729_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11731_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n11733_o = n11731_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11734_o = n11730_o | n11733_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11735_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n11737_o = n11735_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11738_o = n11734_o | n11737_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11739_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n11741_o = n11739_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11742_o = n11738_o | n11741_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11743_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n11745_o = n11743_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11746_o = n11742_o | n11745_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11747_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n11749_o = n11747_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11750_o = n11746_o | n11749_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11751_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n11753_o = n11751_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11754_o = n11750_o | n11753_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n11755_o = ~n11754_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n11756_o = ~n11755_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11768_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n11770_o = n11768_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11772_o = 1'b0 | n11770_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11774_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n11776_o = n11774_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11777_o = n11772_o | n11776_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11778_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n11780_o = n11778_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11781_o = n11777_o | n11780_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11782_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n11784_o = n11782_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11785_o = n11781_o | n11784_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11786_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n11788_o = n11786_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11789_o = n11785_o | n11788_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11790_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n11792_o = n11790_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11793_o = n11789_o | n11792_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11794_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n11796_o = n11794_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11797_o = n11793_o | n11796_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11798_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n11800_o = n11798_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11801_o = n11797_o | n11800_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11802_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n11804_o = n11802_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11805_o = n11801_o | n11804_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11806_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n11808_o = n11806_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11809_o = n11805_o | n11808_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11810_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n11812_o = n11810_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11813_o = n11809_o | n11812_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11814_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n11816_o = n11814_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11817_o = n11813_o | n11816_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11818_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n11820_o = n11818_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11821_o = n11817_o | n11820_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11822_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n11824_o = n11822_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11825_o = n11821_o | n11824_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11826_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n11828_o = n11826_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11829_o = n11825_o | n11828_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11830_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n11832_o = n11830_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11833_o = n11829_o | n11832_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11834_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n11836_o = n11834_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11837_o = n11833_o | n11836_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11838_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n11840_o = n11838_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11841_o = n11837_o | n11840_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11842_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n11844_o = n11842_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11845_o = n11841_o | n11844_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11846_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n11848_o = n11846_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11849_o = n11845_o | n11848_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11850_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n11852_o = n11850_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11853_o = n11849_o | n11852_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11854_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n11856_o = n11854_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11857_o = n11853_o | n11856_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11858_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n11860_o = n11858_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11861_o = n11857_o | n11860_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11862_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n11864_o = n11862_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11865_o = n11861_o | n11864_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11866_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n11868_o = n11866_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11869_o = n11865_o | n11868_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11870_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n11872_o = n11870_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11873_o = n11869_o | n11872_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11874_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n11876_o = n11874_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11877_o = n11873_o | n11876_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11878_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n11880_o = n11878_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11881_o = n11877_o | n11880_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11882_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n11884_o = n11882_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11885_o = n11881_o | n11884_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11886_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n11888_o = n11886_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11889_o = n11885_o | n11888_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11890_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n11892_o = n11890_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11893_o = n11889_o | n11892_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11894_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n11896_o = n11894_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11897_o = n11893_o | n11896_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n11898_o = ~n11897_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n11899_o = ~n11898_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11911_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n11913_o = n11911_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11915_o = 1'b0 | n11913_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11917_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n11919_o = n11917_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11920_o = n11915_o | n11919_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11921_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n11923_o = n11921_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11924_o = n11920_o | n11923_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11925_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n11927_o = n11925_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11928_o = n11924_o | n11927_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11929_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n11931_o = n11929_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11932_o = n11928_o | n11931_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11933_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n11935_o = n11933_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11936_o = n11932_o | n11935_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11937_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n11939_o = n11937_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11940_o = n11936_o | n11939_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11941_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n11943_o = n11941_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11944_o = n11940_o | n11943_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11945_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n11947_o = n11945_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11948_o = n11944_o | n11947_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11949_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n11951_o = n11949_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11952_o = n11948_o | n11951_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11953_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n11955_o = n11953_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n11956_o = n11952_o | n11955_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11957_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n11959_o = n11957_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11960_o = n11956_o | n11959_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11961_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n11963_o = n11961_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11964_o = n11960_o | n11963_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11965_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n11967_o = n11965_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11968_o = n11964_o | n11967_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11969_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n11971_o = n11969_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11972_o = n11968_o | n11971_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11973_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n11975_o = n11973_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11976_o = n11972_o | n11975_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11977_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n11979_o = n11977_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11980_o = n11976_o | n11979_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11981_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n11983_o = n11981_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11984_o = n11980_o | n11983_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11985_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n11987_o = n11985_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11988_o = n11984_o | n11987_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11989_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n11991_o = n11989_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11992_o = n11988_o | n11991_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11993_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n11995_o = n11993_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n11996_o = n11992_o | n11995_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n11997_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n11999_o = n11997_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12000_o = n11996_o | n11999_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12001_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n12003_o = n12001_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12004_o = n12000_o | n12003_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12005_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n12007_o = n12005_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12008_o = n12004_o | n12007_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12009_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n12011_o = n12009_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12012_o = n12008_o | n12011_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12013_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n12015_o = n12013_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12016_o = n12012_o | n12015_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12017_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12019_o = n12017_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12020_o = n12016_o | n12019_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12021_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12023_o = n12021_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12024_o = n12020_o | n12023_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12025_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12027_o = n12025_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12028_o = n12024_o | n12027_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12029_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12031_o = n12029_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12032_o = n12028_o | n12031_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12033_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12035_o = n12033_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12036_o = n12032_o | n12035_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12037_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12039_o = n12037_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12040_o = n12036_o | n12039_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12041_o = ~n12040_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n12042_o = ~n12041_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12054_o = krom_block_rom_block_wl[31];
  /* vlm5030_pack.vhd:50:32  */
  assign n12056_o = n12054_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12058_o = 1'b0 | n12056_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12060_o = krom_block_rom_block_wl[30];
  /* vlm5030_pack.vhd:50:32  */
  assign n12062_o = n12060_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12063_o = n12058_o | n12062_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12064_o = krom_block_rom_block_wl[29];
  /* vlm5030_pack.vhd:50:32  */
  assign n12066_o = n12064_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12067_o = n12063_o | n12066_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12068_o = krom_block_rom_block_wl[28];
  /* vlm5030_pack.vhd:50:32  */
  assign n12070_o = n12068_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12071_o = n12067_o | n12070_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12072_o = krom_block_rom_block_wl[27];
  /* vlm5030_pack.vhd:50:32  */
  assign n12074_o = n12072_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12075_o = n12071_o | n12074_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12076_o = krom_block_rom_block_wl[26];
  /* vlm5030_pack.vhd:50:32  */
  assign n12078_o = n12076_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12079_o = n12075_o | n12078_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12080_o = krom_block_rom_block_wl[25];
  /* vlm5030_pack.vhd:50:32  */
  assign n12082_o = n12080_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12083_o = n12079_o | n12082_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12084_o = krom_block_rom_block_wl[24];
  /* vlm5030_pack.vhd:50:32  */
  assign n12086_o = n12084_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12087_o = n12083_o | n12086_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12088_o = krom_block_rom_block_wl[23];
  /* vlm5030_pack.vhd:50:32  */
  assign n12090_o = n12088_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12091_o = n12087_o | n12090_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12092_o = krom_block_rom_block_wl[22];
  /* vlm5030_pack.vhd:50:32  */
  assign n12094_o = n12092_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12095_o = n12091_o | n12094_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12096_o = krom_block_rom_block_wl[21];
  /* vlm5030_pack.vhd:50:32  */
  assign n12098_o = n12096_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12099_o = n12095_o | n12098_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12100_o = krom_block_rom_block_wl[20];
  /* vlm5030_pack.vhd:50:32  */
  assign n12102_o = n12100_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12103_o = n12099_o | n12102_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12104_o = krom_block_rom_block_wl[19];
  /* vlm5030_pack.vhd:50:32  */
  assign n12106_o = n12104_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12107_o = n12103_o | n12106_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12108_o = krom_block_rom_block_wl[18];
  /* vlm5030_pack.vhd:50:32  */
  assign n12110_o = n12108_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12111_o = n12107_o | n12110_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12112_o = krom_block_rom_block_wl[17];
  /* vlm5030_pack.vhd:50:32  */
  assign n12114_o = n12112_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12115_o = n12111_o | n12114_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12116_o = krom_block_rom_block_wl[16];
  /* vlm5030_pack.vhd:50:32  */
  assign n12118_o = n12116_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12119_o = n12115_o | n12118_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12120_o = krom_block_rom_block_wl[15];
  /* vlm5030_pack.vhd:50:32  */
  assign n12122_o = n12120_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12123_o = n12119_o | n12122_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12124_o = krom_block_rom_block_wl[14];
  /* vlm5030_pack.vhd:50:32  */
  assign n12126_o = n12124_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12127_o = n12123_o | n12126_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12128_o = krom_block_rom_block_wl[13];
  /* vlm5030_pack.vhd:50:32  */
  assign n12130_o = n12128_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12131_o = n12127_o | n12130_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12132_o = krom_block_rom_block_wl[12];
  /* vlm5030_pack.vhd:50:32  */
  assign n12134_o = n12132_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12135_o = n12131_o | n12134_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12136_o = krom_block_rom_block_wl[11];
  /* vlm5030_pack.vhd:50:32  */
  assign n12138_o = n12136_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12139_o = n12135_o | n12138_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12140_o = krom_block_rom_block_wl[10];
  /* vlm5030_pack.vhd:50:32  */
  assign n12142_o = n12140_o & 1'b1;
  /* vlm5030_pack.vhd:50:20  */
  assign n12143_o = n12139_o | n12142_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12144_o = krom_block_rom_block_wl[9];
  /* vlm5030_pack.vhd:50:32  */
  assign n12146_o = n12144_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12147_o = n12143_o | n12146_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12148_o = krom_block_rom_block_wl[8];
  /* vlm5030_pack.vhd:50:32  */
  assign n12150_o = n12148_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12151_o = n12147_o | n12150_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12152_o = krom_block_rom_block_wl[7];
  /* vlm5030_pack.vhd:50:32  */
  assign n12154_o = n12152_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12155_o = n12151_o | n12154_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12156_o = krom_block_rom_block_wl[6];
  /* vlm5030_pack.vhd:50:32  */
  assign n12158_o = n12156_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12159_o = n12155_o | n12158_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12160_o = krom_block_rom_block_wl[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12162_o = n12160_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12163_o = n12159_o | n12162_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12164_o = krom_block_rom_block_wl[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12166_o = n12164_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12167_o = n12163_o | n12166_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12168_o = krom_block_rom_block_wl[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12170_o = n12168_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12171_o = n12167_o | n12170_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12172_o = krom_block_rom_block_wl[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12174_o = n12172_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12175_o = n12171_o | n12174_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12176_o = krom_block_rom_block_wl[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12178_o = n12176_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12179_o = n12175_o | n12178_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12180_o = krom_block_rom_block_wl[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12182_o = n12180_o & 1'b0;
  /* vlm5030_pack.vhd:50:20  */
  assign n12183_o = n12179_o | n12182_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12184_o = ~n12183_o;
  /* vlm5030_pack.vhd:67:12  */
  assign n12185_o = ~n12184_o;
  assign n12189_o = {n12185_o, n12042_o, n11899_o, n11756_o};
  assign n12190_o = {n11613_o, n11470_o, n11327_o, 1'b0};
  assign n12191_o = {1'b0, 1'b0};
  assign n12192_o = {n12189_o, n12190_o, n12191_o};
  /* vlm5030_gl.vhd:1289:21  */
  assign n12193_o = krom_block_ka[1];
  /* vlm5030_gl.vhd:1289:15  */
  assign n12194_o = ~n12193_o;
  /* vlm5030_gl.vhd:1290:21  */
  assign n12195_o = krom_block_ka[2];
  /* vlm5030_gl.vhd:1290:15  */
  assign n12196_o = ~n12195_o;
  /* vlm5030_gl.vhd:1291:21  */
  assign n12197_o = krom_block_ka[3];
  /* vlm5030_gl.vhd:1291:15  */
  assign n12198_o = ~n12197_o;
  /* vlm5030_gl.vhd:1292:21  */
  assign n12199_o = krom_block_ka[4];
  /* vlm5030_gl.vhd:1292:15  */
  assign n12200_o = ~n12199_o;
  assign n12207_o = {n12200_o, n12198_o, n12196_o, n12194_o};
  assign n12208_o = {1'b0, 1'b0, 1'b0, 1'b0};
  assign n12209_o = {1'b0, 1'b0};
  assign n12210_o = {n12207_o, n12208_o, n12209_o};
  /* vlm5030_gl.vhd:1300:31  */
  assign n12212_o = ksa[3:1];
  /* vlm5030_pack.vhd:40:24  */
  assign n12218_o = n12212_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n12220_o = 1'b0 | n12218_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n12222_o = n12212_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n12223_o = n12220_o | n12222_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n12224_o = n12212_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n12225_o = n12223_o | n12224_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n12226_o = ~n12225_o;
  /* vlm5030_gl.vhd:1301:26  */
  assign n12227_o = ksa[2];
  /* vlm5030_gl.vhd:1301:38  */
  assign n12228_o = ksa[3];
  /* vlm5030_gl.vhd:1301:50  */
  assign n12229_o = ksa[1];
  /* vlm5030_gl.vhd:1301:42  */
  assign n12230_o = ~(n12228_o & n12229_o);
  /* vlm5030_gl.vhd:1301:30  */
  assign n12231_o = ~(n12227_o | n12230_o);
  assign n12232_o = dinalq[2];
  /* vlm5030_gl.vhd:1302:23  */
  assign n12233_o = ~n12232_o;
  assign n12234_o = ksa[0];
  /* vlm5030_gl.vhd:1303:23  */
  assign n12235_o = ~n12234_o;
  /* vlm5030_gl.vhd:1319:33  */
  assign n12236_o = krom_block_rom_block_range_s0s1s2 & krom_block_rom_block_nksa0;
  /* vlm5030_gl.vhd:1319:43  */
  assign n12237_o = n12236_o & krom_block_rom_block_nkaodd;
  /* vlm5030_gl.vhd:1320:33  */
  assign n12238_o = krom_block_rom_block_range_s0s1s2 & krom_block_rom_block_nksa0;
  assign n12239_o = dinalq[2];
  /* vlm5030_gl.vhd:1320:43  */
  assign n12240_o = n12238_o & n12239_o;
  /* vlm5030_gl.vhd:1319:55  */
  assign n12241_o = {n12237_o, n12240_o};
  assign n12242_o = ksa[0];
  /* vlm5030_gl.vhd:1321:33  */
  assign n12243_o = krom_block_rom_block_range_s0s1s2 & n12242_o;
  /* vlm5030_gl.vhd:1320:55  */
  assign n12244_o = {n12241_o, n12243_o};
  /* vlm5030_gl.vhd:1322:33  */
  assign n12245_o = krom_block_rom_block_range_s3s4 & krom_block_rom_block_nksa0;
  /* vlm5030_gl.vhd:1321:55  */
  assign n12246_o = {n12244_o, n12245_o};
  assign n12247_o = ksa[0];
  /* vlm5030_gl.vhd:1323:33  */
  assign n12248_o = krom_block_rom_block_range_s3s4 & n12247_o;
  /* vlm5030_gl.vhd:1322:55  */
  assign n12249_o = {n12246_o, n12248_o};
  /* vlm5030_gl.vhd:1324:33  */
  assign n12250_o = ~(krom_block_rom_block_range_s0s1s2 | krom_block_rom_block_range_s3s4);
  /* vlm5030_gl.vhd:1323:55  */
  assign n12251_o = {n12249_o, n12250_o};
  /* vlm5030_gl.vhd:1327:34  */
  assign n12253_o = krom_block_rom_block_kslice0[9];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12254_o = krom_block_rom_block_kslice1[9];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12255_o = {n12253_o, n12254_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12256_o = krom_block_rom_block_kslice2[9];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12257_o = {n12255_o, n12256_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12258_o = krom_block_rom_block_kslice3[9];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12259_o = {n12257_o, n12258_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12260_o = krom_block_rom_block_kslice4[9];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12261_o = {n12259_o, n12260_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12262_o = krom_block_rom_block_kslice5[9];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12263_o = {n12261_o, n12262_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12269_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12270_o = n12263_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12271_o = n12269_o & n12270_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12273_o = 1'b0 | n12271_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12275_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12276_o = n12263_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12277_o = n12275_o & n12276_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12278_o = n12273_o | n12277_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12279_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12280_o = n12263_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12281_o = n12279_o & n12280_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12282_o = n12278_o | n12281_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12283_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12284_o = n12263_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12285_o = n12283_o & n12284_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12286_o = n12282_o | n12285_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12287_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12288_o = n12263_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12289_o = n12287_o & n12288_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12290_o = n12286_o | n12289_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12291_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12292_o = n12263_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12293_o = n12291_o & n12292_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12294_o = n12290_o | n12293_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12295_o = ~n12294_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12297_o = krom_block_rom_block_kslice0[8];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12298_o = krom_block_rom_block_kslice1[8];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12299_o = {n12297_o, n12298_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12300_o = krom_block_rom_block_kslice2[8];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12301_o = {n12299_o, n12300_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12302_o = krom_block_rom_block_kslice3[8];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12303_o = {n12301_o, n12302_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12304_o = krom_block_rom_block_kslice4[8];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12305_o = {n12303_o, n12304_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12306_o = krom_block_rom_block_kslice5[8];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12307_o = {n12305_o, n12306_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12313_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12314_o = n12307_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12315_o = n12313_o & n12314_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12317_o = 1'b0 | n12315_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12319_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12320_o = n12307_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12321_o = n12319_o & n12320_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12322_o = n12317_o | n12321_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12323_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12324_o = n12307_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12325_o = n12323_o & n12324_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12326_o = n12322_o | n12325_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12327_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12328_o = n12307_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12329_o = n12327_o & n12328_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12330_o = n12326_o | n12329_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12331_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12332_o = n12307_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12333_o = n12331_o & n12332_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12334_o = n12330_o | n12333_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12335_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12336_o = n12307_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12337_o = n12335_o & n12336_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12338_o = n12334_o | n12337_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12339_o = ~n12338_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12341_o = krom_block_rom_block_kslice0[7];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12342_o = krom_block_rom_block_kslice1[7];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12343_o = {n12341_o, n12342_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12344_o = krom_block_rom_block_kslice2[7];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12345_o = {n12343_o, n12344_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12346_o = krom_block_rom_block_kslice3[7];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12347_o = {n12345_o, n12346_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12348_o = krom_block_rom_block_kslice4[7];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12349_o = {n12347_o, n12348_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12350_o = krom_block_rom_block_kslice5[7];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12351_o = {n12349_o, n12350_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12357_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12358_o = n12351_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12359_o = n12357_o & n12358_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12361_o = 1'b0 | n12359_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12363_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12364_o = n12351_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12365_o = n12363_o & n12364_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12366_o = n12361_o | n12365_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12367_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12368_o = n12351_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12369_o = n12367_o & n12368_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12370_o = n12366_o | n12369_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12371_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12372_o = n12351_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12373_o = n12371_o & n12372_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12374_o = n12370_o | n12373_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12375_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12376_o = n12351_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12377_o = n12375_o & n12376_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12378_o = n12374_o | n12377_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12379_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12380_o = n12351_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12381_o = n12379_o & n12380_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12382_o = n12378_o | n12381_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12383_o = ~n12382_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12385_o = krom_block_rom_block_kslice0[6];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12386_o = krom_block_rom_block_kslice1[6];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12387_o = {n12385_o, n12386_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12388_o = krom_block_rom_block_kslice2[6];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12389_o = {n12387_o, n12388_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12390_o = krom_block_rom_block_kslice3[6];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12391_o = {n12389_o, n12390_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12392_o = krom_block_rom_block_kslice4[6];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12393_o = {n12391_o, n12392_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12394_o = krom_block_rom_block_kslice5[6];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12395_o = {n12393_o, n12394_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12401_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12402_o = n12395_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12403_o = n12401_o & n12402_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12405_o = 1'b0 | n12403_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12407_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12408_o = n12395_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12409_o = n12407_o & n12408_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12410_o = n12405_o | n12409_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12411_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12412_o = n12395_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12413_o = n12411_o & n12412_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12414_o = n12410_o | n12413_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12415_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12416_o = n12395_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12417_o = n12415_o & n12416_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12418_o = n12414_o | n12417_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12419_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12420_o = n12395_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12421_o = n12419_o & n12420_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12422_o = n12418_o | n12421_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12423_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12424_o = n12395_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12425_o = n12423_o & n12424_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12426_o = n12422_o | n12425_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12427_o = ~n12426_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12429_o = krom_block_rom_block_kslice0[5];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12430_o = krom_block_rom_block_kslice1[5];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12431_o = {n12429_o, n12430_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12432_o = krom_block_rom_block_kslice2[5];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12433_o = {n12431_o, n12432_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12434_o = krom_block_rom_block_kslice3[5];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12435_o = {n12433_o, n12434_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12436_o = krom_block_rom_block_kslice4[5];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12437_o = {n12435_o, n12436_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12438_o = krom_block_rom_block_kslice5[5];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12439_o = {n12437_o, n12438_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12445_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12446_o = n12439_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12447_o = n12445_o & n12446_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12449_o = 1'b0 | n12447_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12451_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12452_o = n12439_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12453_o = n12451_o & n12452_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12454_o = n12449_o | n12453_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12455_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12456_o = n12439_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12457_o = n12455_o & n12456_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12458_o = n12454_o | n12457_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12459_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12460_o = n12439_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12461_o = n12459_o & n12460_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12462_o = n12458_o | n12461_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12463_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12464_o = n12439_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12465_o = n12463_o & n12464_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12466_o = n12462_o | n12465_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12467_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12468_o = n12439_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12469_o = n12467_o & n12468_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12470_o = n12466_o | n12469_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12471_o = ~n12470_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12473_o = krom_block_rom_block_kslice0[4];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12474_o = krom_block_rom_block_kslice1[4];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12475_o = {n12473_o, n12474_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12476_o = krom_block_rom_block_kslice2[4];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12477_o = {n12475_o, n12476_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12478_o = krom_block_rom_block_kslice3[4];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12479_o = {n12477_o, n12478_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12480_o = krom_block_rom_block_kslice4[4];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12481_o = {n12479_o, n12480_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12482_o = krom_block_rom_block_kslice5[4];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12483_o = {n12481_o, n12482_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12489_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12490_o = n12483_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12491_o = n12489_o & n12490_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12493_o = 1'b0 | n12491_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12495_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12496_o = n12483_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12497_o = n12495_o & n12496_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12498_o = n12493_o | n12497_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12499_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12500_o = n12483_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12501_o = n12499_o & n12500_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12502_o = n12498_o | n12501_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12503_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12504_o = n12483_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12505_o = n12503_o & n12504_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12506_o = n12502_o | n12505_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12507_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12508_o = n12483_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12509_o = n12507_o & n12508_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12510_o = n12506_o | n12509_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12511_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12512_o = n12483_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12513_o = n12511_o & n12512_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12514_o = n12510_o | n12513_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12515_o = ~n12514_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12517_o = krom_block_rom_block_kslice0[3];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12518_o = krom_block_rom_block_kslice1[3];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12519_o = {n12517_o, n12518_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12520_o = krom_block_rom_block_kslice2[3];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12521_o = {n12519_o, n12520_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12522_o = krom_block_rom_block_kslice3[3];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12523_o = {n12521_o, n12522_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12524_o = krom_block_rom_block_kslice4[3];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12525_o = {n12523_o, n12524_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12526_o = krom_block_rom_block_kslice5[3];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12527_o = {n12525_o, n12526_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12533_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12534_o = n12527_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12535_o = n12533_o & n12534_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12537_o = 1'b0 | n12535_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12539_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12540_o = n12527_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12541_o = n12539_o & n12540_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12542_o = n12537_o | n12541_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12543_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12544_o = n12527_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12545_o = n12543_o & n12544_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12546_o = n12542_o | n12545_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12547_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12548_o = n12527_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12549_o = n12547_o & n12548_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12550_o = n12546_o | n12549_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12551_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12552_o = n12527_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12553_o = n12551_o & n12552_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12554_o = n12550_o | n12553_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12555_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12556_o = n12527_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12557_o = n12555_o & n12556_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12558_o = n12554_o | n12557_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12559_o = ~n12558_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12561_o = krom_block_rom_block_kslice0[2];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12562_o = krom_block_rom_block_kslice1[2];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12563_o = {n12561_o, n12562_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12564_o = krom_block_rom_block_kslice2[2];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12565_o = {n12563_o, n12564_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12566_o = krom_block_rom_block_kslice3[2];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12567_o = {n12565_o, n12566_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12568_o = krom_block_rom_block_kslice4[2];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12569_o = {n12567_o, n12568_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12570_o = krom_block_rom_block_kslice5[2];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12571_o = {n12569_o, n12570_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12577_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12578_o = n12571_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12579_o = n12577_o & n12578_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12581_o = 1'b0 | n12579_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12583_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12584_o = n12571_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12585_o = n12583_o & n12584_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12586_o = n12581_o | n12585_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12587_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12588_o = n12571_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12589_o = n12587_o & n12588_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12590_o = n12586_o | n12589_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12591_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12592_o = n12571_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12593_o = n12591_o & n12592_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12594_o = n12590_o | n12593_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12595_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12596_o = n12571_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12597_o = n12595_o & n12596_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12598_o = n12594_o | n12597_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12599_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12600_o = n12571_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12601_o = n12599_o & n12600_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12602_o = n12598_o | n12601_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12603_o = ~n12602_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12605_o = krom_block_rom_block_kslice0[1];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12606_o = krom_block_rom_block_kslice1[1];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12607_o = {n12605_o, n12606_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12608_o = krom_block_rom_block_kslice2[1];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12609_o = {n12607_o, n12608_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12610_o = krom_block_rom_block_kslice3[1];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12611_o = {n12609_o, n12610_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12612_o = krom_block_rom_block_kslice4[1];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12613_o = {n12611_o, n12612_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12614_o = krom_block_rom_block_kslice5[1];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12615_o = {n12613_o, n12614_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12621_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12622_o = n12615_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12623_o = n12621_o & n12622_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12625_o = 1'b0 | n12623_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12627_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12628_o = n12615_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12629_o = n12627_o & n12628_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12630_o = n12625_o | n12629_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12631_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12632_o = n12615_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12633_o = n12631_o & n12632_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12634_o = n12630_o | n12633_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12635_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12636_o = n12615_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12637_o = n12635_o & n12636_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12638_o = n12634_o | n12637_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12639_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12640_o = n12615_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12641_o = n12639_o & n12640_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12642_o = n12638_o | n12641_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12643_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12644_o = n12615_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12645_o = n12643_o & n12644_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12646_o = n12642_o | n12645_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12647_o = ~n12646_o;
  /* vlm5030_gl.vhd:1327:34  */
  assign n12649_o = krom_block_rom_block_kslice0[0];
  /* vlm5030_gl.vhd:1328:34  */
  assign n12650_o = krom_block_rom_block_kslice1[0];
  /* vlm5030_gl.vhd:1327:40  */
  assign n12651_o = {n12649_o, n12650_o};
  /* vlm5030_gl.vhd:1329:34  */
  assign n12652_o = krom_block_rom_block_kslice2[0];
  /* vlm5030_gl.vhd:1328:40  */
  assign n12653_o = {n12651_o, n12652_o};
  /* vlm5030_gl.vhd:1330:34  */
  assign n12654_o = krom_block_rom_block_kslice3[0];
  /* vlm5030_gl.vhd:1329:40  */
  assign n12655_o = {n12653_o, n12654_o};
  /* vlm5030_gl.vhd:1331:34  */
  assign n12656_o = krom_block_rom_block_kslice4[0];
  /* vlm5030_gl.vhd:1330:40  */
  assign n12657_o = {n12655_o, n12656_o};
  /* vlm5030_gl.vhd:1332:34  */
  assign n12658_o = krom_block_rom_block_kslice5[0];
  /* vlm5030_gl.vhd:1331:40  */
  assign n12659_o = {n12657_o, n12658_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n12665_o = krom_block_rom_block_wl_slice[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n12666_o = n12659_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n12667_o = n12665_o & n12666_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12669_o = 1'b0 | n12667_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12671_o = krom_block_rom_block_wl_slice[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n12672_o = n12659_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n12673_o = n12671_o & n12672_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12674_o = n12669_o | n12673_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12675_o = krom_block_rom_block_wl_slice[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n12676_o = n12659_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n12677_o = n12675_o & n12676_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12678_o = n12674_o | n12677_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12679_o = krom_block_rom_block_wl_slice[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n12680_o = n12659_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n12681_o = n12679_o & n12680_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12682_o = n12678_o | n12681_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12683_o = krom_block_rom_block_wl_slice[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n12684_o = n12659_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n12685_o = n12683_o & n12684_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12686_o = n12682_o | n12685_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n12687_o = krom_block_rom_block_wl_slice[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n12688_o = n12659_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n12689_o = n12687_o & n12688_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n12690_o = n12686_o | n12689_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n12691_o = ~n12690_o;
  /* vlm5030_gl.vhd:1335:15  */
  assign n12692_o = ~krom_block_rom_block_kout;
  assign n12693_o = {n12295_o, n12339_o, n12383_o, n12427_o, n12471_o, n12515_o, n12559_o, n12603_o, n12647_o, n12691_o};
  /* vlm5030_gl.vhd:1376:12  */
  always @*
    regfile_block_rf0 = n13737_q; // (isignal)
  initial
    regfile_block_rf0 = 10'b0000000000;
  /* vlm5030_gl.vhd:1376:17  */
  always @*
    regfile_block_rf1 = n13739_q; // (isignal)
  initial
    regfile_block_rf1 = 10'b0000000000;
  /* vlm5030_gl.vhd:1377:12  */
  always @*
    regfile_block_rf2 = n13741_q; // (isignal)
  initial
    regfile_block_rf2 = 4'b0000;
  /* vlm5030_gl.vhd:1377:17  */
  always @*
    regfile_block_rf3 = n13743_q; // (isignal)
  initial
    regfile_block_rf3 = 4'b0000;
  /* vlm5030_gl.vhd:1378:12  */
  always @*
    regfile_block_rf4 = n13745_q; // (isignal)
  initial
    regfile_block_rf4 = 3'b000;
  /* vlm5030_gl.vhd:1378:17  */
  always @*
    regfile_block_rf5 = n13747_q; // (isignal)
  initial
    regfile_block_rf5 = 3'b000;
  /* vlm5030_gl.vhd:1379:12  */
  always @*
    regfile_block_rf6 = n13749_q; // (isignal)
  initial
    regfile_block_rf6 = 3'b000;
  /* vlm5030_gl.vhd:1379:17  */
  always @*
    regfile_block_rf7 = n13751_q; // (isignal)
  initial
    regfile_block_rf7 = 3'b000;
  /* vlm5030_gl.vhd:1380:12  */
  always @*
    regfile_block_rf8 = n13753_q; // (isignal)
  initial
    regfile_block_rf8 = 3'b000;
  /* vlm5030_gl.vhd:1380:17  */
  always @*
    regfile_block_rf9 = n13755_q; // (isignal)
  initial
    regfile_block_rf9 = 3'b000;
  /* vlm5030_gl.vhd:1381:12  */
  always @*
    regfile_block_rf10 = n13757_q; // (isignal)
  initial
    regfile_block_rf10 = 7'b0000000;
  /* vlm5030_gl.vhd:1382:12  */
  always @*
    regfile_block_rf11 = n13759_q; // (isignal)
  initial
    regfile_block_rf11 = 7'b0000000;
  /* vlm5030_gl.vhd:1383:12  */
  assign regfile_block_a = n12706_o; // (signal)
  /* vlm5030_gl.vhd:1384:12  */
  assign regfile_block_al = n12796_o; // (signal)
  /* vlm5030_gl.vhd:1385:12  */
  assign regfile_block_nrfdo = n13760_o; // (signal)
  /* vlm5030_gl.vhd:1388:10  */
  assign n12706_o = {26'b0, ksa};  //  uext
  assign n12709_o = osc[0];
  /* vlm5030_gl.vhd:1395:13  */
  assign n12712_o = regfile_block_a == 31'b0000000000000000000000000000000;
  /* vlm5030_gl.vhd:1396:13  */
  assign n12714_o = regfile_block_a == 31'b0000000000000000000000000000001;
  /* vlm5030_gl.vhd:1397:36  */
  assign n12715_o = nkdo[9:6];
  /* vlm5030_gl.vhd:1397:13  */
  assign n12717_o = regfile_block_a == 31'b0000000000000000000000000000010;
  /* vlm5030_gl.vhd:1398:36  */
  assign n12718_o = nkdo[9:6];
  /* vlm5030_gl.vhd:1398:13  */
  assign n12720_o = regfile_block_a == 31'b0000000000000000000000000000011;
  /* vlm5030_gl.vhd:1399:36  */
  assign n12721_o = nkdo[9:7];
  /* vlm5030_gl.vhd:1399:13  */
  assign n12723_o = regfile_block_a == 31'b0000000000000000000000000000100;
  /* vlm5030_gl.vhd:1400:36  */
  assign n12724_o = nkdo[9:7];
  /* vlm5030_gl.vhd:1400:13  */
  assign n12726_o = regfile_block_a == 31'b0000000000000000000000000000101;
  /* vlm5030_gl.vhd:1401:36  */
  assign n12727_o = nkdo[9:7];
  /* vlm5030_gl.vhd:1401:13  */
  assign n12729_o = regfile_block_a == 31'b0000000000000000000000000000110;
  /* vlm5030_gl.vhd:1402:36  */
  assign n12730_o = nkdo[9:7];
  /* vlm5030_gl.vhd:1402:13  */
  assign n12732_o = regfile_block_a == 31'b0000000000000000000000000000111;
  /* vlm5030_gl.vhd:1403:36  */
  assign n12733_o = nkdo[9:7];
  /* vlm5030_gl.vhd:1403:13  */
  assign n12735_o = regfile_block_a == 31'b0000000000000000000000000001000;
  /* vlm5030_gl.vhd:1404:36  */
  assign n12736_o = nkdo[9:7];
  /* vlm5030_gl.vhd:1404:13  */
  assign n12738_o = regfile_block_a == 31'b0000000000000000000000000001001;
  /* vlm5030_gl.vhd:1405:36  */
  assign n12739_o = nkdo[6:0];
  /* vlm5030_gl.vhd:1405:13  */
  assign n12741_o = regfile_block_a == 31'b0000000000000000000000000001010;
  /* vlm5030_gl.vhd:1406:36  */
  assign n12742_o = nkdo[9:3];
  /* vlm5030_gl.vhd:1406:13  */
  assign n12744_o = regfile_block_a == 31'b0000000000000000000000000001011;
  assign n12745_o = {n12744_o, n12741_o, n12738_o, n12735_o, n12732_o, n12729_o, n12726_o, n12723_o, n12720_o, n12717_o, n12714_o, n12712_o};
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12746_o = regfile_block_rf0;
      12'b010000000000: n12746_o = regfile_block_rf0;
      12'b001000000000: n12746_o = regfile_block_rf0;
      12'b000100000000: n12746_o = regfile_block_rf0;
      12'b000010000000: n12746_o = regfile_block_rf0;
      12'b000001000000: n12746_o = regfile_block_rf0;
      12'b000000100000: n12746_o = regfile_block_rf0;
      12'b000000010000: n12746_o = regfile_block_rf0;
      12'b000000001000: n12746_o = regfile_block_rf0;
      12'b000000000100: n12746_o = regfile_block_rf0;
      12'b000000000010: n12746_o = regfile_block_rf0;
      12'b000000000001: n12746_o = nkdo;
      default: n12746_o = regfile_block_rf0;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12747_o = regfile_block_rf1;
      12'b010000000000: n12747_o = regfile_block_rf1;
      12'b001000000000: n12747_o = regfile_block_rf1;
      12'b000100000000: n12747_o = regfile_block_rf1;
      12'b000010000000: n12747_o = regfile_block_rf1;
      12'b000001000000: n12747_o = regfile_block_rf1;
      12'b000000100000: n12747_o = regfile_block_rf1;
      12'b000000010000: n12747_o = regfile_block_rf1;
      12'b000000001000: n12747_o = regfile_block_rf1;
      12'b000000000100: n12747_o = regfile_block_rf1;
      12'b000000000010: n12747_o = nkdo;
      12'b000000000001: n12747_o = regfile_block_rf1;
      default: n12747_o = regfile_block_rf1;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12748_o = regfile_block_rf2;
      12'b010000000000: n12748_o = regfile_block_rf2;
      12'b001000000000: n12748_o = regfile_block_rf2;
      12'b000100000000: n12748_o = regfile_block_rf2;
      12'b000010000000: n12748_o = regfile_block_rf2;
      12'b000001000000: n12748_o = regfile_block_rf2;
      12'b000000100000: n12748_o = regfile_block_rf2;
      12'b000000010000: n12748_o = regfile_block_rf2;
      12'b000000001000: n12748_o = regfile_block_rf2;
      12'b000000000100: n12748_o = n12715_o;
      12'b000000000010: n12748_o = regfile_block_rf2;
      12'b000000000001: n12748_o = regfile_block_rf2;
      default: n12748_o = regfile_block_rf2;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12749_o = regfile_block_rf3;
      12'b010000000000: n12749_o = regfile_block_rf3;
      12'b001000000000: n12749_o = regfile_block_rf3;
      12'b000100000000: n12749_o = regfile_block_rf3;
      12'b000010000000: n12749_o = regfile_block_rf3;
      12'b000001000000: n12749_o = regfile_block_rf3;
      12'b000000100000: n12749_o = regfile_block_rf3;
      12'b000000010000: n12749_o = regfile_block_rf3;
      12'b000000001000: n12749_o = n12718_o;
      12'b000000000100: n12749_o = regfile_block_rf3;
      12'b000000000010: n12749_o = regfile_block_rf3;
      12'b000000000001: n12749_o = regfile_block_rf3;
      default: n12749_o = regfile_block_rf3;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12750_o = regfile_block_rf4;
      12'b010000000000: n12750_o = regfile_block_rf4;
      12'b001000000000: n12750_o = regfile_block_rf4;
      12'b000100000000: n12750_o = regfile_block_rf4;
      12'b000010000000: n12750_o = regfile_block_rf4;
      12'b000001000000: n12750_o = regfile_block_rf4;
      12'b000000100000: n12750_o = regfile_block_rf4;
      12'b000000010000: n12750_o = n12721_o;
      12'b000000001000: n12750_o = regfile_block_rf4;
      12'b000000000100: n12750_o = regfile_block_rf4;
      12'b000000000010: n12750_o = regfile_block_rf4;
      12'b000000000001: n12750_o = regfile_block_rf4;
      default: n12750_o = regfile_block_rf4;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12751_o = regfile_block_rf5;
      12'b010000000000: n12751_o = regfile_block_rf5;
      12'b001000000000: n12751_o = regfile_block_rf5;
      12'b000100000000: n12751_o = regfile_block_rf5;
      12'b000010000000: n12751_o = regfile_block_rf5;
      12'b000001000000: n12751_o = regfile_block_rf5;
      12'b000000100000: n12751_o = n12724_o;
      12'b000000010000: n12751_o = regfile_block_rf5;
      12'b000000001000: n12751_o = regfile_block_rf5;
      12'b000000000100: n12751_o = regfile_block_rf5;
      12'b000000000010: n12751_o = regfile_block_rf5;
      12'b000000000001: n12751_o = regfile_block_rf5;
      default: n12751_o = regfile_block_rf5;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12752_o = regfile_block_rf6;
      12'b010000000000: n12752_o = regfile_block_rf6;
      12'b001000000000: n12752_o = regfile_block_rf6;
      12'b000100000000: n12752_o = regfile_block_rf6;
      12'b000010000000: n12752_o = regfile_block_rf6;
      12'b000001000000: n12752_o = n12727_o;
      12'b000000100000: n12752_o = regfile_block_rf6;
      12'b000000010000: n12752_o = regfile_block_rf6;
      12'b000000001000: n12752_o = regfile_block_rf6;
      12'b000000000100: n12752_o = regfile_block_rf6;
      12'b000000000010: n12752_o = regfile_block_rf6;
      12'b000000000001: n12752_o = regfile_block_rf6;
      default: n12752_o = regfile_block_rf6;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12753_o = regfile_block_rf7;
      12'b010000000000: n12753_o = regfile_block_rf7;
      12'b001000000000: n12753_o = regfile_block_rf7;
      12'b000100000000: n12753_o = regfile_block_rf7;
      12'b000010000000: n12753_o = n12730_o;
      12'b000001000000: n12753_o = regfile_block_rf7;
      12'b000000100000: n12753_o = regfile_block_rf7;
      12'b000000010000: n12753_o = regfile_block_rf7;
      12'b000000001000: n12753_o = regfile_block_rf7;
      12'b000000000100: n12753_o = regfile_block_rf7;
      12'b000000000010: n12753_o = regfile_block_rf7;
      12'b000000000001: n12753_o = regfile_block_rf7;
      default: n12753_o = regfile_block_rf7;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12754_o = regfile_block_rf8;
      12'b010000000000: n12754_o = regfile_block_rf8;
      12'b001000000000: n12754_o = regfile_block_rf8;
      12'b000100000000: n12754_o = n12733_o;
      12'b000010000000: n12754_o = regfile_block_rf8;
      12'b000001000000: n12754_o = regfile_block_rf8;
      12'b000000100000: n12754_o = regfile_block_rf8;
      12'b000000010000: n12754_o = regfile_block_rf8;
      12'b000000001000: n12754_o = regfile_block_rf8;
      12'b000000000100: n12754_o = regfile_block_rf8;
      12'b000000000010: n12754_o = regfile_block_rf8;
      12'b000000000001: n12754_o = regfile_block_rf8;
      default: n12754_o = regfile_block_rf8;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12755_o = regfile_block_rf9;
      12'b010000000000: n12755_o = regfile_block_rf9;
      12'b001000000000: n12755_o = n12736_o;
      12'b000100000000: n12755_o = regfile_block_rf9;
      12'b000010000000: n12755_o = regfile_block_rf9;
      12'b000001000000: n12755_o = regfile_block_rf9;
      12'b000000100000: n12755_o = regfile_block_rf9;
      12'b000000010000: n12755_o = regfile_block_rf9;
      12'b000000001000: n12755_o = regfile_block_rf9;
      12'b000000000100: n12755_o = regfile_block_rf9;
      12'b000000000010: n12755_o = regfile_block_rf9;
      12'b000000000001: n12755_o = regfile_block_rf9;
      default: n12755_o = regfile_block_rf9;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12756_o = regfile_block_rf10;
      12'b010000000000: n12756_o = n12739_o;
      12'b001000000000: n12756_o = regfile_block_rf10;
      12'b000100000000: n12756_o = regfile_block_rf10;
      12'b000010000000: n12756_o = regfile_block_rf10;
      12'b000001000000: n12756_o = regfile_block_rf10;
      12'b000000100000: n12756_o = regfile_block_rf10;
      12'b000000010000: n12756_o = regfile_block_rf10;
      12'b000000001000: n12756_o = regfile_block_rf10;
      12'b000000000100: n12756_o = regfile_block_rf10;
      12'b000000000010: n12756_o = regfile_block_rf10;
      12'b000000000001: n12756_o = regfile_block_rf10;
      default: n12756_o = regfile_block_rf10;
    endcase
  /* vlm5030_gl.vhd:1394:11  */
  always @*
    case (n12745_o)
      12'b100000000000: n12757_o = n12742_o;
      12'b010000000000: n12757_o = regfile_block_rf11;
      12'b001000000000: n12757_o = regfile_block_rf11;
      12'b000100000000: n12757_o = regfile_block_rf11;
      12'b000010000000: n12757_o = regfile_block_rf11;
      12'b000001000000: n12757_o = regfile_block_rf11;
      12'b000000100000: n12757_o = regfile_block_rf11;
      12'b000000010000: n12757_o = regfile_block_rf11;
      12'b000000001000: n12757_o = regfile_block_rf11;
      12'b000000000100: n12757_o = regfile_block_rf11;
      12'b000000000010: n12757_o = regfile_block_rf11;
      12'b000000000001: n12757_o = regfile_block_rf11;
      default: n12757_o = regfile_block_rf11;
    endcase
  /* vlm5030_gl.vhd:1416:12  */
  assign n12785_o = {1'b0, regfile_block_a};  //  uext
  /* vlm5030_gl.vhd:1416:12  */
  assign n12787_o = $signed(n12785_o) <= $signed(32'b00000000000000000000000000001011);
  /* vlm5030_gl.vhd:1417:12  */
  assign n12788_o = regfile_block_a[3:0];  // trunc
  /* vlm5030_gl.vhd:1417:12  */
  assign n12790_o = 4'b1011 - n12788_o;
  /* vlm5030_gl.vhd:1416:7  */
  assign n12796_o = n12787_o ? n20596_o : 12'b000000000000;
  /* vlm5030_gl.vhd:1423:30  */
  assign n12800_o = regfile_block_rf0[0];
  /* vlm5030_gl.vhd:1423:39  */
  assign n12801_o = regfile_block_rf1[0];
  /* vlm5030_gl.vhd:1423:34  */
  assign n12802_o = {n12800_o, n12801_o};
  /* vlm5030_gl.vhd:1423:43  */
  assign n12804_o = {n12802_o, 1'b1};
  /* vlm5030_gl.vhd:1423:52  */
  assign n12806_o = {n12804_o, 1'b1};
  /* vlm5030_gl.vhd:1423:61  */
  assign n12808_o = {n12806_o, 1'b1};
  /* vlm5030_gl.vhd:1423:70  */
  assign n12810_o = {n12808_o, 1'b1};
  /* vlm5030_gl.vhd:1423:79  */
  assign n12812_o = {n12810_o, 1'b1};
  /* vlm5030_gl.vhd:1423:88  */
  assign n12814_o = {n12812_o, 1'b1};
  /* vlm5030_gl.vhd:1423:97  */
  assign n12816_o = {n12814_o, 1'b1};
  /* vlm5030_gl.vhd:1423:106  */
  assign n12818_o = {n12816_o, 1'b1};
  /* vlm5030_gl.vhd:1423:121  */
  assign n12819_o = regfile_block_rf10[0];
  /* vlm5030_gl.vhd:1423:115  */
  assign n12820_o = {n12818_o, n12819_o};
  /* vlm5030_gl.vhd:1423:125  */
  assign n12822_o = {n12820_o, 1'b1};
  /* vlm5030_pack.vhd:60:26  */
  assign n12828_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n12829_o = n12822_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n12830_o = ~n12829_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12831_o = n12828_o & n12830_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12833_o = 1'b0 | n12831_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12835_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n12836_o = n12822_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n12837_o = ~n12836_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12838_o = n12835_o & n12837_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12839_o = n12833_o | n12838_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12840_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n12841_o = n12822_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n12842_o = ~n12841_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12843_o = n12840_o & n12842_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12844_o = n12839_o | n12843_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12845_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n12846_o = n12822_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n12847_o = ~n12846_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12848_o = n12845_o & n12847_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12849_o = n12844_o | n12848_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12850_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n12851_o = n12822_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n12852_o = ~n12851_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12853_o = n12850_o & n12852_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12854_o = n12849_o | n12853_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12855_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n12856_o = n12822_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n12857_o = ~n12856_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12858_o = n12855_o & n12857_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12859_o = n12854_o | n12858_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12860_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n12861_o = n12822_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n12862_o = ~n12861_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12863_o = n12860_o & n12862_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12864_o = n12859_o | n12863_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12865_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n12866_o = n12822_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n12867_o = ~n12866_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12868_o = n12865_o & n12867_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12869_o = n12864_o | n12868_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12870_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n12871_o = n12822_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n12872_o = ~n12871_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12873_o = n12870_o & n12872_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12874_o = n12869_o | n12873_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12875_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n12876_o = n12822_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n12877_o = ~n12876_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12878_o = n12875_o & n12877_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12879_o = n12874_o | n12878_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12880_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n12881_o = n12822_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n12882_o = ~n12881_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12883_o = n12880_o & n12882_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12884_o = n12879_o | n12883_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12885_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n12886_o = n12822_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n12887_o = ~n12886_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12888_o = n12885_o & n12887_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12889_o = n12884_o | n12888_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n12890_o = ~n12889_o;
  /* vlm5030_gl.vhd:1424:30  */
  assign n12892_o = regfile_block_rf0[1];
  /* vlm5030_gl.vhd:1424:39  */
  assign n12893_o = regfile_block_rf1[1];
  /* vlm5030_gl.vhd:1424:34  */
  assign n12894_o = {n12892_o, n12893_o};
  /* vlm5030_gl.vhd:1424:43  */
  assign n12896_o = {n12894_o, 1'b1};
  /* vlm5030_gl.vhd:1424:52  */
  assign n12898_o = {n12896_o, 1'b1};
  /* vlm5030_gl.vhd:1424:61  */
  assign n12900_o = {n12898_o, 1'b1};
  /* vlm5030_gl.vhd:1424:70  */
  assign n12902_o = {n12900_o, 1'b1};
  /* vlm5030_gl.vhd:1424:79  */
  assign n12904_o = {n12902_o, 1'b1};
  /* vlm5030_gl.vhd:1424:88  */
  assign n12906_o = {n12904_o, 1'b1};
  /* vlm5030_gl.vhd:1424:97  */
  assign n12908_o = {n12906_o, 1'b1};
  /* vlm5030_gl.vhd:1424:106  */
  assign n12910_o = {n12908_o, 1'b1};
  /* vlm5030_gl.vhd:1424:121  */
  assign n12911_o = regfile_block_rf10[1];
  /* vlm5030_gl.vhd:1424:115  */
  assign n12912_o = {n12910_o, n12911_o};
  /* vlm5030_gl.vhd:1424:125  */
  assign n12914_o = {n12912_o, 1'b1};
  /* vlm5030_pack.vhd:60:26  */
  assign n12920_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n12921_o = n12914_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n12922_o = ~n12921_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12923_o = n12920_o & n12922_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12925_o = 1'b0 | n12923_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12927_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n12928_o = n12914_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n12929_o = ~n12928_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12930_o = n12927_o & n12929_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12931_o = n12925_o | n12930_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12932_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n12933_o = n12914_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n12934_o = ~n12933_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12935_o = n12932_o & n12934_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12936_o = n12931_o | n12935_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12937_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n12938_o = n12914_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n12939_o = ~n12938_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12940_o = n12937_o & n12939_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12941_o = n12936_o | n12940_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12942_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n12943_o = n12914_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n12944_o = ~n12943_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12945_o = n12942_o & n12944_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12946_o = n12941_o | n12945_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12947_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n12948_o = n12914_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n12949_o = ~n12948_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12950_o = n12947_o & n12949_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12951_o = n12946_o | n12950_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12952_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n12953_o = n12914_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n12954_o = ~n12953_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12955_o = n12952_o & n12954_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12956_o = n12951_o | n12955_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12957_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n12958_o = n12914_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n12959_o = ~n12958_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12960_o = n12957_o & n12959_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12961_o = n12956_o | n12960_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12962_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n12963_o = n12914_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n12964_o = ~n12963_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12965_o = n12962_o & n12964_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12966_o = n12961_o | n12965_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12967_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n12968_o = n12914_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n12969_o = ~n12968_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12970_o = n12967_o & n12969_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12971_o = n12966_o | n12970_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12972_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n12973_o = n12914_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n12974_o = ~n12973_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12975_o = n12972_o & n12974_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12976_o = n12971_o | n12975_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n12977_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n12978_o = n12914_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n12979_o = ~n12978_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n12980_o = n12977_o & n12979_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n12981_o = n12976_o | n12980_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n12982_o = ~n12981_o;
  /* vlm5030_gl.vhd:1425:30  */
  assign n12984_o = regfile_block_rf0[2];
  /* vlm5030_gl.vhd:1425:39  */
  assign n12985_o = regfile_block_rf1[2];
  /* vlm5030_gl.vhd:1425:34  */
  assign n12986_o = {n12984_o, n12985_o};
  /* vlm5030_gl.vhd:1425:43  */
  assign n12988_o = {n12986_o, 1'b1};
  /* vlm5030_gl.vhd:1425:52  */
  assign n12990_o = {n12988_o, 1'b1};
  /* vlm5030_gl.vhd:1425:61  */
  assign n12992_o = {n12990_o, 1'b1};
  /* vlm5030_gl.vhd:1425:70  */
  assign n12994_o = {n12992_o, 1'b1};
  /* vlm5030_gl.vhd:1425:79  */
  assign n12996_o = {n12994_o, 1'b1};
  /* vlm5030_gl.vhd:1425:88  */
  assign n12998_o = {n12996_o, 1'b1};
  /* vlm5030_gl.vhd:1425:97  */
  assign n13000_o = {n12998_o, 1'b1};
  /* vlm5030_gl.vhd:1425:106  */
  assign n13002_o = {n13000_o, 1'b1};
  /* vlm5030_gl.vhd:1425:121  */
  assign n13003_o = regfile_block_rf10[2];
  /* vlm5030_gl.vhd:1425:115  */
  assign n13004_o = {n13002_o, n13003_o};
  /* vlm5030_gl.vhd:1425:125  */
  assign n13006_o = {n13004_o, 1'b1};
  /* vlm5030_pack.vhd:60:26  */
  assign n13012_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n13013_o = n13006_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n13014_o = ~n13013_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13015_o = n13012_o & n13014_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13017_o = 1'b0 | n13015_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13019_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n13020_o = n13006_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n13021_o = ~n13020_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13022_o = n13019_o & n13021_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13023_o = n13017_o | n13022_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13024_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n13025_o = n13006_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n13026_o = ~n13025_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13027_o = n13024_o & n13026_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13028_o = n13023_o | n13027_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13029_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n13030_o = n13006_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n13031_o = ~n13030_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13032_o = n13029_o & n13031_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13033_o = n13028_o | n13032_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13034_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n13035_o = n13006_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n13036_o = ~n13035_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13037_o = n13034_o & n13036_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13038_o = n13033_o | n13037_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13039_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n13040_o = n13006_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n13041_o = ~n13040_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13042_o = n13039_o & n13041_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13043_o = n13038_o | n13042_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13044_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n13045_o = n13006_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n13046_o = ~n13045_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13047_o = n13044_o & n13046_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13048_o = n13043_o | n13047_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13049_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n13050_o = n13006_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n13051_o = ~n13050_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13052_o = n13049_o & n13051_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13053_o = n13048_o | n13052_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13054_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n13055_o = n13006_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n13056_o = ~n13055_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13057_o = n13054_o & n13056_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13058_o = n13053_o | n13057_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13059_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n13060_o = n13006_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n13061_o = ~n13060_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13062_o = n13059_o & n13061_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13063_o = n13058_o | n13062_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13064_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n13065_o = n13006_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n13066_o = ~n13065_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13067_o = n13064_o & n13066_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13068_o = n13063_o | n13067_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13069_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n13070_o = n13006_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n13071_o = ~n13070_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13072_o = n13069_o & n13071_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13073_o = n13068_o | n13072_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n13074_o = ~n13073_o;
  /* vlm5030_gl.vhd:1426:30  */
  assign n13076_o = regfile_block_rf0[3];
  /* vlm5030_gl.vhd:1426:39  */
  assign n13077_o = regfile_block_rf1[3];
  /* vlm5030_gl.vhd:1426:34  */
  assign n13078_o = {n13076_o, n13077_o};
  /* vlm5030_gl.vhd:1426:43  */
  assign n13080_o = {n13078_o, 1'b1};
  /* vlm5030_gl.vhd:1426:52  */
  assign n13082_o = {n13080_o, 1'b1};
  /* vlm5030_gl.vhd:1426:61  */
  assign n13084_o = {n13082_o, 1'b1};
  /* vlm5030_gl.vhd:1426:70  */
  assign n13086_o = {n13084_o, 1'b1};
  /* vlm5030_gl.vhd:1426:79  */
  assign n13088_o = {n13086_o, 1'b1};
  /* vlm5030_gl.vhd:1426:88  */
  assign n13090_o = {n13088_o, 1'b1};
  /* vlm5030_gl.vhd:1426:97  */
  assign n13092_o = {n13090_o, 1'b1};
  /* vlm5030_gl.vhd:1426:106  */
  assign n13094_o = {n13092_o, 1'b1};
  /* vlm5030_gl.vhd:1426:121  */
  assign n13095_o = regfile_block_rf10[3];
  /* vlm5030_gl.vhd:1426:115  */
  assign n13096_o = {n13094_o, n13095_o};
  /* vlm5030_gl.vhd:1426:131  */
  assign n13097_o = regfile_block_rf11[0];
  /* vlm5030_gl.vhd:1426:125  */
  assign n13098_o = {n13096_o, n13097_o};
  /* vlm5030_pack.vhd:60:26  */
  assign n13104_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n13105_o = n13098_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n13106_o = ~n13105_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13107_o = n13104_o & n13106_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13109_o = 1'b0 | n13107_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13111_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n13112_o = n13098_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n13113_o = ~n13112_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13114_o = n13111_o & n13113_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13115_o = n13109_o | n13114_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13116_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n13117_o = n13098_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n13118_o = ~n13117_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13119_o = n13116_o & n13118_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13120_o = n13115_o | n13119_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13121_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n13122_o = n13098_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n13123_o = ~n13122_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13124_o = n13121_o & n13123_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13125_o = n13120_o | n13124_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13126_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n13127_o = n13098_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n13128_o = ~n13127_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13129_o = n13126_o & n13128_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13130_o = n13125_o | n13129_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13131_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n13132_o = n13098_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n13133_o = ~n13132_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13134_o = n13131_o & n13133_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13135_o = n13130_o | n13134_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13136_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n13137_o = n13098_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n13138_o = ~n13137_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13139_o = n13136_o & n13138_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13140_o = n13135_o | n13139_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13141_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n13142_o = n13098_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n13143_o = ~n13142_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13144_o = n13141_o & n13143_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13145_o = n13140_o | n13144_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13146_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n13147_o = n13098_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n13148_o = ~n13147_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13149_o = n13146_o & n13148_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13150_o = n13145_o | n13149_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13151_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n13152_o = n13098_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n13153_o = ~n13152_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13154_o = n13151_o & n13153_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13155_o = n13150_o | n13154_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13156_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n13157_o = n13098_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n13158_o = ~n13157_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13159_o = n13156_o & n13158_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13160_o = n13155_o | n13159_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13161_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n13162_o = n13098_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n13163_o = ~n13162_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13164_o = n13161_o & n13163_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13165_o = n13160_o | n13164_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n13166_o = ~n13165_o;
  /* vlm5030_gl.vhd:1427:30  */
  assign n13168_o = regfile_block_rf0[4];
  /* vlm5030_gl.vhd:1427:39  */
  assign n13169_o = regfile_block_rf1[4];
  /* vlm5030_gl.vhd:1427:34  */
  assign n13170_o = {n13168_o, n13169_o};
  /* vlm5030_gl.vhd:1427:43  */
  assign n13172_o = {n13170_o, 1'b1};
  /* vlm5030_gl.vhd:1427:52  */
  assign n13174_o = {n13172_o, 1'b1};
  /* vlm5030_gl.vhd:1427:61  */
  assign n13176_o = {n13174_o, 1'b1};
  /* vlm5030_gl.vhd:1427:70  */
  assign n13178_o = {n13176_o, 1'b1};
  /* vlm5030_gl.vhd:1427:79  */
  assign n13180_o = {n13178_o, 1'b1};
  /* vlm5030_gl.vhd:1427:88  */
  assign n13182_o = {n13180_o, 1'b1};
  /* vlm5030_gl.vhd:1427:97  */
  assign n13184_o = {n13182_o, 1'b1};
  /* vlm5030_gl.vhd:1427:106  */
  assign n13186_o = {n13184_o, 1'b1};
  /* vlm5030_gl.vhd:1427:121  */
  assign n13187_o = regfile_block_rf10[4];
  /* vlm5030_gl.vhd:1427:115  */
  assign n13188_o = {n13186_o, n13187_o};
  /* vlm5030_gl.vhd:1427:131  */
  assign n13189_o = regfile_block_rf11[1];
  /* vlm5030_gl.vhd:1427:125  */
  assign n13190_o = {n13188_o, n13189_o};
  /* vlm5030_pack.vhd:60:26  */
  assign n13196_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n13197_o = n13190_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n13198_o = ~n13197_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13199_o = n13196_o & n13198_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13201_o = 1'b0 | n13199_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13203_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n13204_o = n13190_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n13205_o = ~n13204_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13206_o = n13203_o & n13205_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13207_o = n13201_o | n13206_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13208_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n13209_o = n13190_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n13210_o = ~n13209_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13211_o = n13208_o & n13210_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13212_o = n13207_o | n13211_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13213_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n13214_o = n13190_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n13215_o = ~n13214_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13216_o = n13213_o & n13215_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13217_o = n13212_o | n13216_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13218_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n13219_o = n13190_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n13220_o = ~n13219_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13221_o = n13218_o & n13220_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13222_o = n13217_o | n13221_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13223_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n13224_o = n13190_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n13225_o = ~n13224_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13226_o = n13223_o & n13225_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13227_o = n13222_o | n13226_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13228_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n13229_o = n13190_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n13230_o = ~n13229_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13231_o = n13228_o & n13230_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13232_o = n13227_o | n13231_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13233_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n13234_o = n13190_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n13235_o = ~n13234_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13236_o = n13233_o & n13235_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13237_o = n13232_o | n13236_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13238_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n13239_o = n13190_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n13240_o = ~n13239_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13241_o = n13238_o & n13240_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13242_o = n13237_o | n13241_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13243_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n13244_o = n13190_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n13245_o = ~n13244_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13246_o = n13243_o & n13245_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13247_o = n13242_o | n13246_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13248_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n13249_o = n13190_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n13250_o = ~n13249_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13251_o = n13248_o & n13250_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13252_o = n13247_o | n13251_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13253_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n13254_o = n13190_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n13255_o = ~n13254_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13256_o = n13253_o & n13255_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13257_o = n13252_o | n13256_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n13258_o = ~n13257_o;
  /* vlm5030_gl.vhd:1428:30  */
  assign n13260_o = regfile_block_rf0[5];
  /* vlm5030_gl.vhd:1428:39  */
  assign n13261_o = regfile_block_rf1[5];
  /* vlm5030_gl.vhd:1428:34  */
  assign n13262_o = {n13260_o, n13261_o};
  /* vlm5030_gl.vhd:1428:43  */
  assign n13264_o = {n13262_o, 1'b1};
  /* vlm5030_gl.vhd:1428:52  */
  assign n13266_o = {n13264_o, 1'b1};
  /* vlm5030_gl.vhd:1428:61  */
  assign n13268_o = {n13266_o, 1'b1};
  /* vlm5030_gl.vhd:1428:70  */
  assign n13270_o = {n13268_o, 1'b1};
  /* vlm5030_gl.vhd:1428:79  */
  assign n13272_o = {n13270_o, 1'b1};
  /* vlm5030_gl.vhd:1428:88  */
  assign n13274_o = {n13272_o, 1'b1};
  /* vlm5030_gl.vhd:1428:97  */
  assign n13276_o = {n13274_o, 1'b1};
  /* vlm5030_gl.vhd:1428:106  */
  assign n13278_o = {n13276_o, 1'b1};
  /* vlm5030_gl.vhd:1428:121  */
  assign n13279_o = regfile_block_rf10[5];
  /* vlm5030_gl.vhd:1428:115  */
  assign n13280_o = {n13278_o, n13279_o};
  /* vlm5030_gl.vhd:1428:131  */
  assign n13281_o = regfile_block_rf11[2];
  /* vlm5030_gl.vhd:1428:125  */
  assign n13282_o = {n13280_o, n13281_o};
  /* vlm5030_pack.vhd:60:26  */
  assign n13288_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n13289_o = n13282_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n13290_o = ~n13289_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13291_o = n13288_o & n13290_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13293_o = 1'b0 | n13291_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13295_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n13296_o = n13282_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n13297_o = ~n13296_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13298_o = n13295_o & n13297_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13299_o = n13293_o | n13298_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13300_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n13301_o = n13282_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n13302_o = ~n13301_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13303_o = n13300_o & n13302_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13304_o = n13299_o | n13303_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13305_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n13306_o = n13282_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n13307_o = ~n13306_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13308_o = n13305_o & n13307_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13309_o = n13304_o | n13308_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13310_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n13311_o = n13282_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n13312_o = ~n13311_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13313_o = n13310_o & n13312_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13314_o = n13309_o | n13313_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13315_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n13316_o = n13282_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n13317_o = ~n13316_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13318_o = n13315_o & n13317_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13319_o = n13314_o | n13318_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13320_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n13321_o = n13282_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n13322_o = ~n13321_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13323_o = n13320_o & n13322_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13324_o = n13319_o | n13323_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13325_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n13326_o = n13282_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n13327_o = ~n13326_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13328_o = n13325_o & n13327_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13329_o = n13324_o | n13328_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13330_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n13331_o = n13282_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n13332_o = ~n13331_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13333_o = n13330_o & n13332_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13334_o = n13329_o | n13333_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13335_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n13336_o = n13282_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n13337_o = ~n13336_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13338_o = n13335_o & n13337_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13339_o = n13334_o | n13338_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13340_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n13341_o = n13282_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n13342_o = ~n13341_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13343_o = n13340_o & n13342_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13344_o = n13339_o | n13343_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13345_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n13346_o = n13282_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n13347_o = ~n13346_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13348_o = n13345_o & n13347_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13349_o = n13344_o | n13348_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n13350_o = ~n13349_o;
  /* vlm5030_gl.vhd:1429:30  */
  assign n13352_o = regfile_block_rf0[6];
  /* vlm5030_gl.vhd:1429:39  */
  assign n13353_o = regfile_block_rf1[6];
  /* vlm5030_gl.vhd:1429:34  */
  assign n13354_o = {n13352_o, n13353_o};
  /* vlm5030_gl.vhd:1429:48  */
  assign n13355_o = regfile_block_rf2[0];
  /* vlm5030_gl.vhd:1429:43  */
  assign n13356_o = {n13354_o, n13355_o};
  /* vlm5030_gl.vhd:1429:57  */
  assign n13357_o = regfile_block_rf3[0];
  /* vlm5030_gl.vhd:1429:52  */
  assign n13358_o = {n13356_o, n13357_o};
  /* vlm5030_gl.vhd:1429:61  */
  assign n13360_o = {n13358_o, 1'b1};
  /* vlm5030_gl.vhd:1429:70  */
  assign n13362_o = {n13360_o, 1'b1};
  /* vlm5030_gl.vhd:1429:79  */
  assign n13364_o = {n13362_o, 1'b1};
  /* vlm5030_gl.vhd:1429:88  */
  assign n13366_o = {n13364_o, 1'b1};
  /* vlm5030_gl.vhd:1429:97  */
  assign n13368_o = {n13366_o, 1'b1};
  /* vlm5030_gl.vhd:1429:106  */
  assign n13370_o = {n13368_o, 1'b1};
  /* vlm5030_gl.vhd:1429:121  */
  assign n13371_o = regfile_block_rf10[6];
  /* vlm5030_gl.vhd:1429:115  */
  assign n13372_o = {n13370_o, n13371_o};
  /* vlm5030_gl.vhd:1429:131  */
  assign n13373_o = regfile_block_rf11[3];
  /* vlm5030_gl.vhd:1429:125  */
  assign n13374_o = {n13372_o, n13373_o};
  /* vlm5030_pack.vhd:60:26  */
  assign n13380_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n13381_o = n13374_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n13382_o = ~n13381_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13383_o = n13380_o & n13382_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13385_o = 1'b0 | n13383_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13387_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n13388_o = n13374_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n13389_o = ~n13388_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13390_o = n13387_o & n13389_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13391_o = n13385_o | n13390_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13392_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n13393_o = n13374_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n13394_o = ~n13393_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13395_o = n13392_o & n13394_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13396_o = n13391_o | n13395_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13397_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n13398_o = n13374_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n13399_o = ~n13398_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13400_o = n13397_o & n13399_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13401_o = n13396_o | n13400_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13402_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n13403_o = n13374_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n13404_o = ~n13403_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13405_o = n13402_o & n13404_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13406_o = n13401_o | n13405_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13407_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n13408_o = n13374_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n13409_o = ~n13408_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13410_o = n13407_o & n13409_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13411_o = n13406_o | n13410_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13412_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n13413_o = n13374_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n13414_o = ~n13413_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13415_o = n13412_o & n13414_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13416_o = n13411_o | n13415_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13417_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n13418_o = n13374_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n13419_o = ~n13418_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13420_o = n13417_o & n13419_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13421_o = n13416_o | n13420_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13422_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n13423_o = n13374_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n13424_o = ~n13423_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13425_o = n13422_o & n13424_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13426_o = n13421_o | n13425_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13427_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n13428_o = n13374_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n13429_o = ~n13428_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13430_o = n13427_o & n13429_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13431_o = n13426_o | n13430_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13432_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n13433_o = n13374_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n13434_o = ~n13433_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13435_o = n13432_o & n13434_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13436_o = n13431_o | n13435_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13437_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n13438_o = n13374_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n13439_o = ~n13438_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13440_o = n13437_o & n13439_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13441_o = n13436_o | n13440_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n13442_o = ~n13441_o;
  /* vlm5030_gl.vhd:1430:30  */
  assign n13444_o = regfile_block_rf0[7];
  /* vlm5030_gl.vhd:1430:39  */
  assign n13445_o = regfile_block_rf1[7];
  /* vlm5030_gl.vhd:1430:34  */
  assign n13446_o = {n13444_o, n13445_o};
  /* vlm5030_gl.vhd:1430:48  */
  assign n13447_o = regfile_block_rf2[1];
  /* vlm5030_gl.vhd:1430:43  */
  assign n13448_o = {n13446_o, n13447_o};
  /* vlm5030_gl.vhd:1430:57  */
  assign n13449_o = regfile_block_rf3[1];
  /* vlm5030_gl.vhd:1430:52  */
  assign n13450_o = {n13448_o, n13449_o};
  /* vlm5030_gl.vhd:1430:66  */
  assign n13451_o = regfile_block_rf4[0];
  /* vlm5030_gl.vhd:1430:61  */
  assign n13452_o = {n13450_o, n13451_o};
  /* vlm5030_gl.vhd:1430:75  */
  assign n13453_o = regfile_block_rf5[0];
  /* vlm5030_gl.vhd:1430:70  */
  assign n13454_o = {n13452_o, n13453_o};
  /* vlm5030_gl.vhd:1430:84  */
  assign n13455_o = regfile_block_rf6[0];
  /* vlm5030_gl.vhd:1430:79  */
  assign n13456_o = {n13454_o, n13455_o};
  /* vlm5030_gl.vhd:1430:93  */
  assign n13457_o = regfile_block_rf7[0];
  /* vlm5030_gl.vhd:1430:88  */
  assign n13458_o = {n13456_o, n13457_o};
  /* vlm5030_gl.vhd:1430:102  */
  assign n13459_o = regfile_block_rf8[0];
  /* vlm5030_gl.vhd:1430:97  */
  assign n13460_o = {n13458_o, n13459_o};
  /* vlm5030_gl.vhd:1430:111  */
  assign n13461_o = regfile_block_rf9[0];
  /* vlm5030_gl.vhd:1430:106  */
  assign n13462_o = {n13460_o, n13461_o};
  /* vlm5030_gl.vhd:1430:115  */
  assign n13464_o = {n13462_o, 1'b1};
  /* vlm5030_gl.vhd:1430:131  */
  assign n13465_o = regfile_block_rf11[4];
  /* vlm5030_gl.vhd:1430:125  */
  assign n13466_o = {n13464_o, n13465_o};
  /* vlm5030_pack.vhd:60:26  */
  assign n13472_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n13473_o = n13466_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n13474_o = ~n13473_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13475_o = n13472_o & n13474_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13477_o = 1'b0 | n13475_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13479_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n13480_o = n13466_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n13481_o = ~n13480_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13482_o = n13479_o & n13481_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13483_o = n13477_o | n13482_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13484_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n13485_o = n13466_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n13486_o = ~n13485_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13487_o = n13484_o & n13486_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13488_o = n13483_o | n13487_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13489_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n13490_o = n13466_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n13491_o = ~n13490_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13492_o = n13489_o & n13491_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13493_o = n13488_o | n13492_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13494_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n13495_o = n13466_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n13496_o = ~n13495_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13497_o = n13494_o & n13496_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13498_o = n13493_o | n13497_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13499_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n13500_o = n13466_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n13501_o = ~n13500_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13502_o = n13499_o & n13501_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13503_o = n13498_o | n13502_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13504_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n13505_o = n13466_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n13506_o = ~n13505_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13507_o = n13504_o & n13506_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13508_o = n13503_o | n13507_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13509_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n13510_o = n13466_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n13511_o = ~n13510_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13512_o = n13509_o & n13511_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13513_o = n13508_o | n13512_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13514_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n13515_o = n13466_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n13516_o = ~n13515_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13517_o = n13514_o & n13516_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13518_o = n13513_o | n13517_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13519_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n13520_o = n13466_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n13521_o = ~n13520_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13522_o = n13519_o & n13521_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13523_o = n13518_o | n13522_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13524_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n13525_o = n13466_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n13526_o = ~n13525_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13527_o = n13524_o & n13526_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13528_o = n13523_o | n13527_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13529_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n13530_o = n13466_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n13531_o = ~n13530_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13532_o = n13529_o & n13531_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13533_o = n13528_o | n13532_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n13534_o = ~n13533_o;
  /* vlm5030_gl.vhd:1431:30  */
  assign n13536_o = regfile_block_rf0[8];
  /* vlm5030_gl.vhd:1431:39  */
  assign n13537_o = regfile_block_rf1[8];
  /* vlm5030_gl.vhd:1431:34  */
  assign n13538_o = {n13536_o, n13537_o};
  /* vlm5030_gl.vhd:1431:48  */
  assign n13539_o = regfile_block_rf2[2];
  /* vlm5030_gl.vhd:1431:43  */
  assign n13540_o = {n13538_o, n13539_o};
  /* vlm5030_gl.vhd:1431:57  */
  assign n13541_o = regfile_block_rf3[2];
  /* vlm5030_gl.vhd:1431:52  */
  assign n13542_o = {n13540_o, n13541_o};
  /* vlm5030_gl.vhd:1431:66  */
  assign n13543_o = regfile_block_rf4[1];
  /* vlm5030_gl.vhd:1431:61  */
  assign n13544_o = {n13542_o, n13543_o};
  /* vlm5030_gl.vhd:1431:75  */
  assign n13545_o = regfile_block_rf5[1];
  /* vlm5030_gl.vhd:1431:70  */
  assign n13546_o = {n13544_o, n13545_o};
  /* vlm5030_gl.vhd:1431:84  */
  assign n13547_o = regfile_block_rf6[1];
  /* vlm5030_gl.vhd:1431:79  */
  assign n13548_o = {n13546_o, n13547_o};
  /* vlm5030_gl.vhd:1431:93  */
  assign n13549_o = regfile_block_rf7[1];
  /* vlm5030_gl.vhd:1431:88  */
  assign n13550_o = {n13548_o, n13549_o};
  /* vlm5030_gl.vhd:1431:102  */
  assign n13551_o = regfile_block_rf8[1];
  /* vlm5030_gl.vhd:1431:97  */
  assign n13552_o = {n13550_o, n13551_o};
  /* vlm5030_gl.vhd:1431:111  */
  assign n13553_o = regfile_block_rf9[1];
  /* vlm5030_gl.vhd:1431:106  */
  assign n13554_o = {n13552_o, n13553_o};
  /* vlm5030_gl.vhd:1431:115  */
  assign n13556_o = {n13554_o, 1'b1};
  /* vlm5030_gl.vhd:1431:131  */
  assign n13557_o = regfile_block_rf11[5];
  /* vlm5030_gl.vhd:1431:125  */
  assign n13558_o = {n13556_o, n13557_o};
  /* vlm5030_pack.vhd:60:26  */
  assign n13564_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n13565_o = n13558_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n13566_o = ~n13565_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13567_o = n13564_o & n13566_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13569_o = 1'b0 | n13567_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13571_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n13572_o = n13558_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n13573_o = ~n13572_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13574_o = n13571_o & n13573_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13575_o = n13569_o | n13574_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13576_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n13577_o = n13558_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n13578_o = ~n13577_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13579_o = n13576_o & n13578_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13580_o = n13575_o | n13579_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13581_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n13582_o = n13558_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n13583_o = ~n13582_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13584_o = n13581_o & n13583_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13585_o = n13580_o | n13584_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13586_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n13587_o = n13558_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n13588_o = ~n13587_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13589_o = n13586_o & n13588_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13590_o = n13585_o | n13589_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13591_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n13592_o = n13558_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n13593_o = ~n13592_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13594_o = n13591_o & n13593_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13595_o = n13590_o | n13594_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13596_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n13597_o = n13558_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n13598_o = ~n13597_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13599_o = n13596_o & n13598_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13600_o = n13595_o | n13599_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13601_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n13602_o = n13558_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n13603_o = ~n13602_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13604_o = n13601_o & n13603_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13605_o = n13600_o | n13604_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13606_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n13607_o = n13558_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n13608_o = ~n13607_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13609_o = n13606_o & n13608_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13610_o = n13605_o | n13609_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13611_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n13612_o = n13558_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n13613_o = ~n13612_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13614_o = n13611_o & n13613_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13615_o = n13610_o | n13614_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13616_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n13617_o = n13558_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n13618_o = ~n13617_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13619_o = n13616_o & n13618_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13620_o = n13615_o | n13619_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13621_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n13622_o = n13558_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n13623_o = ~n13622_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13624_o = n13621_o & n13623_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13625_o = n13620_o | n13624_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n13626_o = ~n13625_o;
  /* vlm5030_gl.vhd:1432:30  */
  assign n13628_o = regfile_block_rf0[9];
  /* vlm5030_gl.vhd:1432:39  */
  assign n13629_o = regfile_block_rf1[9];
  /* vlm5030_gl.vhd:1432:34  */
  assign n13630_o = {n13628_o, n13629_o};
  /* vlm5030_gl.vhd:1432:48  */
  assign n13631_o = regfile_block_rf2[3];
  /* vlm5030_gl.vhd:1432:43  */
  assign n13632_o = {n13630_o, n13631_o};
  /* vlm5030_gl.vhd:1432:57  */
  assign n13633_o = regfile_block_rf3[3];
  /* vlm5030_gl.vhd:1432:52  */
  assign n13634_o = {n13632_o, n13633_o};
  /* vlm5030_gl.vhd:1432:66  */
  assign n13635_o = regfile_block_rf4[2];
  /* vlm5030_gl.vhd:1432:61  */
  assign n13636_o = {n13634_o, n13635_o};
  /* vlm5030_gl.vhd:1432:75  */
  assign n13637_o = regfile_block_rf5[2];
  /* vlm5030_gl.vhd:1432:70  */
  assign n13638_o = {n13636_o, n13637_o};
  /* vlm5030_gl.vhd:1432:84  */
  assign n13639_o = regfile_block_rf6[2];
  /* vlm5030_gl.vhd:1432:79  */
  assign n13640_o = {n13638_o, n13639_o};
  /* vlm5030_gl.vhd:1432:93  */
  assign n13641_o = regfile_block_rf7[2];
  /* vlm5030_gl.vhd:1432:88  */
  assign n13642_o = {n13640_o, n13641_o};
  /* vlm5030_gl.vhd:1432:102  */
  assign n13643_o = regfile_block_rf8[2];
  /* vlm5030_gl.vhd:1432:97  */
  assign n13644_o = {n13642_o, n13643_o};
  /* vlm5030_gl.vhd:1432:111  */
  assign n13645_o = regfile_block_rf9[2];
  /* vlm5030_gl.vhd:1432:106  */
  assign n13646_o = {n13644_o, n13645_o};
  /* vlm5030_gl.vhd:1432:115  */
  assign n13648_o = {n13646_o, 1'b1};
  /* vlm5030_gl.vhd:1432:131  */
  assign n13649_o = regfile_block_rf11[6];
  /* vlm5030_gl.vhd:1432:125  */
  assign n13650_o = {n13648_o, n13649_o};
  /* vlm5030_pack.vhd:60:26  */
  assign n13656_o = regfile_block_al[11];
  /* vlm5030_pack.vhd:60:43  */
  assign n13657_o = n13650_o[11];
  /* vlm5030_pack.vhd:60:36  */
  assign n13658_o = ~n13657_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13659_o = n13656_o & n13658_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13661_o = 1'b0 | n13659_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13663_o = regfile_block_al[10];
  /* vlm5030_pack.vhd:60:43  */
  assign n13664_o = n13650_o[10];
  /* vlm5030_pack.vhd:60:36  */
  assign n13665_o = ~n13664_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13666_o = n13663_o & n13665_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13667_o = n13661_o | n13666_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13668_o = regfile_block_al[9];
  /* vlm5030_pack.vhd:60:43  */
  assign n13669_o = n13650_o[9];
  /* vlm5030_pack.vhd:60:36  */
  assign n13670_o = ~n13669_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13671_o = n13668_o & n13670_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13672_o = n13667_o | n13671_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13673_o = regfile_block_al[8];
  /* vlm5030_pack.vhd:60:43  */
  assign n13674_o = n13650_o[8];
  /* vlm5030_pack.vhd:60:36  */
  assign n13675_o = ~n13674_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13676_o = n13673_o & n13675_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13677_o = n13672_o | n13676_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13678_o = regfile_block_al[7];
  /* vlm5030_pack.vhd:60:43  */
  assign n13679_o = n13650_o[7];
  /* vlm5030_pack.vhd:60:36  */
  assign n13680_o = ~n13679_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13681_o = n13678_o & n13680_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13682_o = n13677_o | n13681_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13683_o = regfile_block_al[6];
  /* vlm5030_pack.vhd:60:43  */
  assign n13684_o = n13650_o[6];
  /* vlm5030_pack.vhd:60:36  */
  assign n13685_o = ~n13684_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13686_o = n13683_o & n13685_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13687_o = n13682_o | n13686_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13688_o = regfile_block_al[5];
  /* vlm5030_pack.vhd:60:43  */
  assign n13689_o = n13650_o[5];
  /* vlm5030_pack.vhd:60:36  */
  assign n13690_o = ~n13689_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13691_o = n13688_o & n13690_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13692_o = n13687_o | n13691_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13693_o = regfile_block_al[4];
  /* vlm5030_pack.vhd:60:43  */
  assign n13694_o = n13650_o[4];
  /* vlm5030_pack.vhd:60:36  */
  assign n13695_o = ~n13694_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13696_o = n13693_o & n13695_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13697_o = n13692_o | n13696_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13698_o = regfile_block_al[3];
  /* vlm5030_pack.vhd:60:43  */
  assign n13699_o = n13650_o[3];
  /* vlm5030_pack.vhd:60:36  */
  assign n13700_o = ~n13699_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13701_o = n13698_o & n13700_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13702_o = n13697_o | n13701_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13703_o = regfile_block_al[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n13704_o = n13650_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n13705_o = ~n13704_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13706_o = n13703_o & n13705_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13707_o = n13702_o | n13706_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13708_o = regfile_block_al[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n13709_o = n13650_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n13710_o = ~n13709_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13711_o = n13708_o & n13710_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13712_o = n13707_o | n13711_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n13713_o = regfile_block_al[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n13714_o = n13650_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n13715_o = ~n13714_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n13716_o = n13713_o & n13715_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n13717_o = n13712_o | n13716_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n13718_o = ~n13717_o;
  /* vlm5030_gl.vhd:1434:13  */
  assign n13719_o = ~regfile_block_nrfdo;
  /* vlm5030_gl.vhd:1436:28  */
  assign n13721_o = rfdo[9:7];
  /* vlm5030_pack.vhd:40:24  */
  assign n13727_o = n13721_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n13729_o = 1'b0 | n13727_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n13731_o = n13721_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n13732_o = n13729_o | n13731_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n13733_o = n13721_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n13734_o = n13732_o | n13733_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n13735_o = ~n13734_o;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13736_o = rflatchwen ? n12746_o : regfile_block_rf0;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13737_q <= n13736_o;
  initial
    n13737_q = 10'b0000000000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13738_o = rflatchwen ? n12747_o : regfile_block_rf1;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13739_q <= n13738_o;
  initial
    n13739_q = 10'b0000000000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13740_o = rflatchwen ? n12748_o : regfile_block_rf2;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13741_q <= n13740_o;
  initial
    n13741_q = 4'b0000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13742_o = rflatchwen ? n12749_o : regfile_block_rf3;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13743_q <= n13742_o;
  initial
    n13743_q = 4'b0000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13744_o = rflatchwen ? n12750_o : regfile_block_rf4;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13745_q <= n13744_o;
  initial
    n13745_q = 3'b000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13746_o = rflatchwen ? n12751_o : regfile_block_rf5;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13747_q <= n13746_o;
  initial
    n13747_q = 3'b000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13748_o = rflatchwen ? n12752_o : regfile_block_rf6;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13749_q <= n13748_o;
  initial
    n13749_q = 3'b000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13750_o = rflatchwen ? n12753_o : regfile_block_rf7;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13751_q <= n13750_o;
  initial
    n13751_q = 3'b000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13752_o = rflatchwen ? n12754_o : regfile_block_rf8;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13753_q <= n13752_o;
  initial
    n13753_q = 3'b000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13754_o = rflatchwen ? n12755_o : regfile_block_rf9;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13755_q <= n13754_o;
  initial
    n13755_q = 3'b000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13756_o = rflatchwen ? n12756_o : regfile_block_rf10;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13757_q <= n13756_o;
  initial
    n13757_q = 7'b0000000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13758_o = rflatchwen ? n12757_o : regfile_block_rf11;
  /* vlm5030_gl.vhd:1392:7  */
  always @(posedge n12709_o)
    n13759_q <= n13758_o;
  initial
    n13759_q = 7'b0000000;
  /* vlm5030_gl.vhd:1392:7  */
  assign n13760_o = {n13718_o, n13626_o, n13534_o, n13442_o, n13350_o, n13258_o, n13166_o, n13074_o, n12982_o, n12890_o};
  /* vlm5030_gl.vhd:1446:12  */
  assign addshift_block_nidlat = n14455_o; // (signal)
  /* vlm5030_gl.vhd:1446:20  */
  assign addshift_block_port_nid = n14456_o; // (signal)
  /* vlm5030_gl.vhd:1447:12  */
  assign addshift_block_port_rf = n14457_o; // (signal)
  /* vlm5030_gl.vhd:1448:12  */
  assign addshift_block_sumlat = n14491_o; // (signal)
  /* vlm5030_gl.vhd:1449:12  */
  assign addshift_block_cin = n14492_o; // (signal)
  /* vlm5030_gl.vhd:1449:17  */
  assign addshift_block_sum = n14493_o; // (signal)
  /* vlm5030_gl.vhd:1450:12  */
  assign addshift_block_idpos = n13770_o; // (signal)
  /* vlm5030_gl.vhd:1453:22  */
  assign n13762_o = dq[6];
  /* vlm5030_gl.vhd:1453:26  */
  assign n13763_o = n13762_o & updtpitch;
  /* clock_functions_pack.vhd:170:25  */
  assign n13768_o = c2d5fin[1];
  /* clock_functions_pack.vhd:170:16  */
  assign n13769_o = ~(n13763_o | n13768_o);
  /* vlm5030_gl.vhd:1453:14  */
  assign n13770_o = ~n13769_o;
  /* vlm5030_gl.vhd:1455:15  */
  assign n13771_o = ~addshift_block_idpos;
  assign n13774_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n13781_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n13782_o = nid[9];
  /* vlm5030_gl.vhd:1473:34  */
  assign n13788_o = addshift_block_nidlat[9];
  /* vlm5030_gl.vhd:1473:24  */
  assign n13789_o = ~n13788_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n13790_o = addshift_block_idpos ? n13789_o : n13791_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n13791_o = addshift_block_nidlat[9];
  /* vlm5030_gl.vhd:1475:28  */
  assign n13792_o = rfdo[9];
  /* clock_functions_pack.vhd:175:17  */
  assign n13798_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n13799_o = ~n13798_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n13800_o = n13799_o ? n13792_o : n13803_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n13801_o = addshift_block_sumlat[10];
  /* vlm5030_gl.vhd:1476:52  */
  assign n13802_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n13803_o = n13802_o ? n13801_o : n13804_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n13804_o = addshift_block_sumlat[11];
  /* vlm5030_gl.vhd:1479:29  */
  assign n13805_o = addshift_block_port_nid[9];
  /* vlm5030_gl.vhd:1479:46  */
  assign n13806_o = addshift_block_port_rf[9];
  /* vlm5030_gl.vhd:1479:35  */
  assign n13807_o = n13805_o ^ n13806_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n13808_o = addshift_block_cin[9];
  /* vlm5030_gl.vhd:1479:52  */
  assign n13809_o = n13807_o ^ n13808_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n13810_o = addshift_block_port_nid[9];
  /* vlm5030_gl.vhd:1481:47  */
  assign n13811_o = addshift_block_port_rf[9];
  /* vlm5030_gl.vhd:1481:36  */
  assign n13812_o = n13810_o & n13811_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n13813_o = addshift_block_port_nid[9];
  /* vlm5030_gl.vhd:1481:83  */
  assign n13814_o = addshift_block_port_rf[9];
  /* vlm5030_gl.vhd:1481:73  */
  assign n13815_o = n13813_o | n13814_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n13816_o = addshift_block_cin[9];
  /* vlm5030_gl.vhd:1481:90  */
  assign n13817_o = n13815_o & n13816_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n13818_o = n13812_o | n13817_o;
  assign n13821_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n13828_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n13829_o = addshift_block_sum[9];
  assign n13837_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n13844_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n13845_o = nid[8];
  /* vlm5030_gl.vhd:1473:34  */
  assign n13851_o = addshift_block_nidlat[8];
  /* vlm5030_gl.vhd:1473:24  */
  assign n13852_o = ~n13851_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n13853_o = addshift_block_idpos ? n13852_o : n13854_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n13854_o = addshift_block_nidlat[8];
  /* vlm5030_gl.vhd:1475:28  */
  assign n13855_o = rfdo[8];
  /* clock_functions_pack.vhd:175:17  */
  assign n13861_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n13862_o = ~n13861_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n13863_o = n13862_o ? n13855_o : n13866_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n13864_o = addshift_block_sumlat[9];
  /* vlm5030_gl.vhd:1476:52  */
  assign n13865_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n13866_o = n13865_o ? n13864_o : n13867_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n13867_o = addshift_block_sumlat[10];
  /* vlm5030_gl.vhd:1479:29  */
  assign n13868_o = addshift_block_port_nid[8];
  /* vlm5030_gl.vhd:1479:46  */
  assign n13869_o = addshift_block_port_rf[8];
  /* vlm5030_gl.vhd:1479:35  */
  assign n13870_o = n13868_o ^ n13869_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n13871_o = addshift_block_cin[8];
  /* vlm5030_gl.vhd:1479:52  */
  assign n13872_o = n13870_o ^ n13871_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n13873_o = addshift_block_port_nid[8];
  /* vlm5030_gl.vhd:1481:47  */
  assign n13874_o = addshift_block_port_rf[8];
  /* vlm5030_gl.vhd:1481:36  */
  assign n13875_o = n13873_o & n13874_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n13876_o = addshift_block_port_nid[8];
  /* vlm5030_gl.vhd:1481:83  */
  assign n13877_o = addshift_block_port_rf[8];
  /* vlm5030_gl.vhd:1481:73  */
  assign n13878_o = n13876_o | n13877_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n13879_o = addshift_block_cin[8];
  /* vlm5030_gl.vhd:1481:90  */
  assign n13880_o = n13878_o & n13879_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n13881_o = n13875_o | n13880_o;
  assign n13884_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n13891_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n13892_o = addshift_block_sum[8];
  assign n13900_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n13907_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n13908_o = nid[7];
  /* vlm5030_gl.vhd:1473:34  */
  assign n13914_o = addshift_block_nidlat[7];
  /* vlm5030_gl.vhd:1473:24  */
  assign n13915_o = ~n13914_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n13916_o = addshift_block_idpos ? n13915_o : n13917_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n13917_o = addshift_block_nidlat[7];
  /* vlm5030_gl.vhd:1475:28  */
  assign n13918_o = rfdo[7];
  /* clock_functions_pack.vhd:175:17  */
  assign n13924_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n13925_o = ~n13924_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n13926_o = n13925_o ? n13918_o : n13929_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n13927_o = addshift_block_sumlat[8];
  /* vlm5030_gl.vhd:1476:52  */
  assign n13928_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n13929_o = n13928_o ? n13927_o : n13930_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n13930_o = addshift_block_sumlat[9];
  /* vlm5030_gl.vhd:1479:29  */
  assign n13931_o = addshift_block_port_nid[7];
  /* vlm5030_gl.vhd:1479:46  */
  assign n13932_o = addshift_block_port_rf[7];
  /* vlm5030_gl.vhd:1479:35  */
  assign n13933_o = n13931_o ^ n13932_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n13934_o = addshift_block_cin[7];
  /* vlm5030_gl.vhd:1479:52  */
  assign n13935_o = n13933_o ^ n13934_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n13936_o = addshift_block_port_nid[7];
  /* vlm5030_gl.vhd:1481:47  */
  assign n13937_o = addshift_block_port_rf[7];
  /* vlm5030_gl.vhd:1481:36  */
  assign n13938_o = n13936_o & n13937_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n13939_o = addshift_block_port_nid[7];
  /* vlm5030_gl.vhd:1481:83  */
  assign n13940_o = addshift_block_port_rf[7];
  /* vlm5030_gl.vhd:1481:73  */
  assign n13941_o = n13939_o | n13940_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n13942_o = addshift_block_cin[7];
  /* vlm5030_gl.vhd:1481:90  */
  assign n13943_o = n13941_o & n13942_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n13944_o = n13938_o | n13943_o;
  assign n13947_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n13954_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n13955_o = addshift_block_sum[7];
  assign n13963_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n13970_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n13971_o = nid[6];
  /* vlm5030_gl.vhd:1473:34  */
  assign n13977_o = addshift_block_nidlat[6];
  /* vlm5030_gl.vhd:1473:24  */
  assign n13978_o = ~n13977_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n13979_o = addshift_block_idpos ? n13978_o : n13980_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n13980_o = addshift_block_nidlat[6];
  /* vlm5030_gl.vhd:1475:28  */
  assign n13981_o = rfdo[6];
  /* clock_functions_pack.vhd:175:17  */
  assign n13987_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n13988_o = ~n13987_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n13989_o = n13988_o ? n13981_o : n13992_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n13990_o = addshift_block_sumlat[7];
  /* vlm5030_gl.vhd:1476:52  */
  assign n13991_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n13992_o = n13991_o ? n13990_o : n13993_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n13993_o = addshift_block_sumlat[8];
  /* vlm5030_gl.vhd:1479:29  */
  assign n13994_o = addshift_block_port_nid[6];
  /* vlm5030_gl.vhd:1479:46  */
  assign n13995_o = addshift_block_port_rf[6];
  /* vlm5030_gl.vhd:1479:35  */
  assign n13996_o = n13994_o ^ n13995_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n13997_o = addshift_block_cin[6];
  /* vlm5030_gl.vhd:1479:52  */
  assign n13998_o = n13996_o ^ n13997_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n13999_o = addshift_block_port_nid[6];
  /* vlm5030_gl.vhd:1481:47  */
  assign n14000_o = addshift_block_port_rf[6];
  /* vlm5030_gl.vhd:1481:36  */
  assign n14001_o = n13999_o & n14000_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n14002_o = addshift_block_port_nid[6];
  /* vlm5030_gl.vhd:1481:83  */
  assign n14003_o = addshift_block_port_rf[6];
  /* vlm5030_gl.vhd:1481:73  */
  assign n14004_o = n14002_o | n14003_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n14005_o = addshift_block_cin[6];
  /* vlm5030_gl.vhd:1481:90  */
  assign n14006_o = n14004_o & n14005_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n14007_o = n14001_o | n14006_o;
  assign n14010_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14017_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n14018_o = addshift_block_sum[6];
  assign n14026_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14033_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n14034_o = nid[5];
  /* vlm5030_gl.vhd:1473:34  */
  assign n14040_o = addshift_block_nidlat[5];
  /* vlm5030_gl.vhd:1473:24  */
  assign n14041_o = ~n14040_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n14042_o = addshift_block_idpos ? n14041_o : n14043_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n14043_o = addshift_block_nidlat[5];
  /* vlm5030_gl.vhd:1475:28  */
  assign n14044_o = rfdo[5];
  /* clock_functions_pack.vhd:175:17  */
  assign n14050_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n14051_o = ~n14050_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n14052_o = n14051_o ? n14044_o : n14055_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n14053_o = addshift_block_sumlat[6];
  /* vlm5030_gl.vhd:1476:52  */
  assign n14054_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n14055_o = n14054_o ? n14053_o : n14056_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n14056_o = addshift_block_sumlat[7];
  /* vlm5030_gl.vhd:1479:29  */
  assign n14057_o = addshift_block_port_nid[5];
  /* vlm5030_gl.vhd:1479:46  */
  assign n14058_o = addshift_block_port_rf[5];
  /* vlm5030_gl.vhd:1479:35  */
  assign n14059_o = n14057_o ^ n14058_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n14060_o = addshift_block_cin[5];
  /* vlm5030_gl.vhd:1479:52  */
  assign n14061_o = n14059_o ^ n14060_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n14062_o = addshift_block_port_nid[5];
  /* vlm5030_gl.vhd:1481:47  */
  assign n14063_o = addshift_block_port_rf[5];
  /* vlm5030_gl.vhd:1481:36  */
  assign n14064_o = n14062_o & n14063_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n14065_o = addshift_block_port_nid[5];
  /* vlm5030_gl.vhd:1481:83  */
  assign n14066_o = addshift_block_port_rf[5];
  /* vlm5030_gl.vhd:1481:73  */
  assign n14067_o = n14065_o | n14066_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n14068_o = addshift_block_cin[5];
  /* vlm5030_gl.vhd:1481:90  */
  assign n14069_o = n14067_o & n14068_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n14070_o = n14064_o | n14069_o;
  assign n14073_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14080_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n14081_o = addshift_block_sum[5];
  assign n14089_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14096_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n14097_o = nid[4];
  /* vlm5030_gl.vhd:1473:34  */
  assign n14103_o = addshift_block_nidlat[4];
  /* vlm5030_gl.vhd:1473:24  */
  assign n14104_o = ~n14103_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n14105_o = addshift_block_idpos ? n14104_o : n14106_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n14106_o = addshift_block_nidlat[4];
  /* vlm5030_gl.vhd:1475:28  */
  assign n14107_o = rfdo[4];
  /* clock_functions_pack.vhd:175:17  */
  assign n14113_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n14114_o = ~n14113_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n14115_o = n14114_o ? n14107_o : n14118_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n14116_o = addshift_block_sumlat[5];
  /* vlm5030_gl.vhd:1476:52  */
  assign n14117_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n14118_o = n14117_o ? n14116_o : n14119_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n14119_o = addshift_block_sumlat[6];
  /* vlm5030_gl.vhd:1479:29  */
  assign n14120_o = addshift_block_port_nid[4];
  /* vlm5030_gl.vhd:1479:46  */
  assign n14121_o = addshift_block_port_rf[4];
  /* vlm5030_gl.vhd:1479:35  */
  assign n14122_o = n14120_o ^ n14121_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n14123_o = addshift_block_cin[4];
  /* vlm5030_gl.vhd:1479:52  */
  assign n14124_o = n14122_o ^ n14123_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n14125_o = addshift_block_port_nid[4];
  /* vlm5030_gl.vhd:1481:47  */
  assign n14126_o = addshift_block_port_rf[4];
  /* vlm5030_gl.vhd:1481:36  */
  assign n14127_o = n14125_o & n14126_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n14128_o = addshift_block_port_nid[4];
  /* vlm5030_gl.vhd:1481:83  */
  assign n14129_o = addshift_block_port_rf[4];
  /* vlm5030_gl.vhd:1481:73  */
  assign n14130_o = n14128_o | n14129_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n14131_o = addshift_block_cin[4];
  /* vlm5030_gl.vhd:1481:90  */
  assign n14132_o = n14130_o & n14131_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n14133_o = n14127_o | n14132_o;
  assign n14136_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14143_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n14144_o = addshift_block_sum[4];
  assign n14152_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14159_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n14160_o = nid[3];
  /* vlm5030_gl.vhd:1473:34  */
  assign n14166_o = addshift_block_nidlat[3];
  /* vlm5030_gl.vhd:1473:24  */
  assign n14167_o = ~n14166_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n14168_o = addshift_block_idpos ? n14167_o : n14169_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n14169_o = addshift_block_nidlat[3];
  /* vlm5030_gl.vhd:1475:28  */
  assign n14170_o = rfdo[3];
  /* clock_functions_pack.vhd:175:17  */
  assign n14176_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n14177_o = ~n14176_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n14178_o = n14177_o ? n14170_o : n14181_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n14179_o = addshift_block_sumlat[4];
  /* vlm5030_gl.vhd:1476:52  */
  assign n14180_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n14181_o = n14180_o ? n14179_o : n14182_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n14182_o = addshift_block_sumlat[5];
  /* vlm5030_gl.vhd:1479:29  */
  assign n14183_o = addshift_block_port_nid[3];
  /* vlm5030_gl.vhd:1479:46  */
  assign n14184_o = addshift_block_port_rf[3];
  /* vlm5030_gl.vhd:1479:35  */
  assign n14185_o = n14183_o ^ n14184_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n14186_o = addshift_block_cin[3];
  /* vlm5030_gl.vhd:1479:52  */
  assign n14187_o = n14185_o ^ n14186_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n14188_o = addshift_block_port_nid[3];
  /* vlm5030_gl.vhd:1481:47  */
  assign n14189_o = addshift_block_port_rf[3];
  /* vlm5030_gl.vhd:1481:36  */
  assign n14190_o = n14188_o & n14189_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n14191_o = addshift_block_port_nid[3];
  /* vlm5030_gl.vhd:1481:83  */
  assign n14192_o = addshift_block_port_rf[3];
  /* vlm5030_gl.vhd:1481:73  */
  assign n14193_o = n14191_o | n14192_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n14194_o = addshift_block_cin[3];
  /* vlm5030_gl.vhd:1481:90  */
  assign n14195_o = n14193_o & n14194_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n14196_o = n14190_o | n14195_o;
  assign n14199_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14206_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n14207_o = addshift_block_sum[3];
  assign n14215_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14222_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n14223_o = nid[2];
  /* vlm5030_gl.vhd:1473:34  */
  assign n14229_o = addshift_block_nidlat[2];
  /* vlm5030_gl.vhd:1473:24  */
  assign n14230_o = ~n14229_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n14231_o = addshift_block_idpos ? n14230_o : n14232_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n14232_o = addshift_block_nidlat[2];
  /* vlm5030_gl.vhd:1475:28  */
  assign n14233_o = rfdo[2];
  /* clock_functions_pack.vhd:175:17  */
  assign n14239_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n14240_o = ~n14239_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n14241_o = n14240_o ? n14233_o : n14244_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n14242_o = addshift_block_sumlat[3];
  /* vlm5030_gl.vhd:1476:52  */
  assign n14243_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n14244_o = n14243_o ? n14242_o : n14245_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n14245_o = addshift_block_sumlat[4];
  /* vlm5030_gl.vhd:1479:29  */
  assign n14246_o = addshift_block_port_nid[2];
  /* vlm5030_gl.vhd:1479:46  */
  assign n14247_o = addshift_block_port_rf[2];
  /* vlm5030_gl.vhd:1479:35  */
  assign n14248_o = n14246_o ^ n14247_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n14249_o = addshift_block_cin[2];
  /* vlm5030_gl.vhd:1479:52  */
  assign n14250_o = n14248_o ^ n14249_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n14251_o = addshift_block_port_nid[2];
  /* vlm5030_gl.vhd:1481:47  */
  assign n14252_o = addshift_block_port_rf[2];
  /* vlm5030_gl.vhd:1481:36  */
  assign n14253_o = n14251_o & n14252_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n14254_o = addshift_block_port_nid[2];
  /* vlm5030_gl.vhd:1481:83  */
  assign n14255_o = addshift_block_port_rf[2];
  /* vlm5030_gl.vhd:1481:73  */
  assign n14256_o = n14254_o | n14255_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n14257_o = addshift_block_cin[2];
  /* vlm5030_gl.vhd:1481:90  */
  assign n14258_o = n14256_o & n14257_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n14259_o = n14253_o | n14258_o;
  assign n14262_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14269_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n14270_o = addshift_block_sum[2];
  assign n14278_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14285_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n14286_o = nid[1];
  /* vlm5030_gl.vhd:1473:34  */
  assign n14292_o = addshift_block_nidlat[1];
  /* vlm5030_gl.vhd:1473:24  */
  assign n14293_o = ~n14292_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n14294_o = addshift_block_idpos ? n14293_o : n14295_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n14295_o = addshift_block_nidlat[1];
  /* vlm5030_gl.vhd:1475:28  */
  assign n14296_o = rfdo[1];
  /* clock_functions_pack.vhd:175:17  */
  assign n14302_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n14303_o = ~n14302_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n14304_o = n14303_o ? n14296_o : n14307_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n14305_o = addshift_block_sumlat[2];
  /* vlm5030_gl.vhd:1476:52  */
  assign n14306_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n14307_o = n14306_o ? n14305_o : n14308_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n14308_o = addshift_block_sumlat[3];
  /* vlm5030_gl.vhd:1479:29  */
  assign n14309_o = addshift_block_port_nid[1];
  /* vlm5030_gl.vhd:1479:46  */
  assign n14310_o = addshift_block_port_rf[1];
  /* vlm5030_gl.vhd:1479:35  */
  assign n14311_o = n14309_o ^ n14310_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n14312_o = addshift_block_cin[1];
  /* vlm5030_gl.vhd:1479:52  */
  assign n14313_o = n14311_o ^ n14312_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n14314_o = addshift_block_port_nid[1];
  /* vlm5030_gl.vhd:1481:47  */
  assign n14315_o = addshift_block_port_rf[1];
  /* vlm5030_gl.vhd:1481:36  */
  assign n14316_o = n14314_o & n14315_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n14317_o = addshift_block_port_nid[1];
  /* vlm5030_gl.vhd:1481:83  */
  assign n14318_o = addshift_block_port_rf[1];
  /* vlm5030_gl.vhd:1481:73  */
  assign n14319_o = n14317_o | n14318_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n14320_o = addshift_block_cin[1];
  /* vlm5030_gl.vhd:1481:90  */
  assign n14321_o = n14319_o & n14320_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n14322_o = n14316_o | n14321_o;
  assign n14325_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14332_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n14333_o = addshift_block_sum[1];
  assign n14341_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14348_o = c2d1[1];
  /* vlm5030_gl.vhd:1467:31  */
  assign n14349_o = nid[0];
  /* vlm5030_gl.vhd:1473:34  */
  assign n14355_o = addshift_block_nidlat[0];
  /* vlm5030_gl.vhd:1473:24  */
  assign n14356_o = ~n14355_o;
  /* vlm5030_gl.vhd:1473:40  */
  assign n14357_o = addshift_block_idpos ? n14356_o : n14358_o;
  /* vlm5030_gl.vhd:1473:68  */
  assign n14358_o = addshift_block_nidlat[0];
  /* vlm5030_gl.vhd:1475:28  */
  assign n14359_o = rfdo[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14365_o = c2d5fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n14366_o = ~n14365_o;
  /* vlm5030_gl.vhd:1475:38  */
  assign n14367_o = n14366_o ? n14359_o : n14370_o;
  /* vlm5030_gl.vhd:1476:30  */
  assign n14368_o = addshift_block_sumlat[1];
  /* vlm5030_gl.vhd:1476:52  */
  assign n14369_o = ~asshift2;
  /* vlm5030_gl.vhd:1475:58  */
  assign n14370_o = n14369_o ? n14368_o : n14371_o;
  /* vlm5030_gl.vhd:1477:30  */
  assign n14371_o = addshift_block_sumlat[2];
  /* vlm5030_gl.vhd:1479:29  */
  assign n14372_o = addshift_block_port_nid[0];
  /* vlm5030_gl.vhd:1479:46  */
  assign n14373_o = addshift_block_port_rf[0];
  /* vlm5030_gl.vhd:1479:35  */
  assign n14374_o = n14372_o ^ n14373_o;
  /* vlm5030_gl.vhd:1479:59  */
  assign n14375_o = addshift_block_cin[0];
  /* vlm5030_gl.vhd:1479:52  */
  assign n14376_o = n14374_o ^ n14375_o;
  /* vlm5030_gl.vhd:1481:30  */
  assign n14377_o = addshift_block_port_nid[0];
  /* vlm5030_gl.vhd:1481:47  */
  assign n14378_o = addshift_block_port_rf[0];
  /* vlm5030_gl.vhd:1481:36  */
  assign n14379_o = n14377_o & n14378_o;
  /* vlm5030_gl.vhd:1481:67  */
  assign n14380_o = addshift_block_port_nid[0];
  /* vlm5030_gl.vhd:1481:83  */
  assign n14381_o = addshift_block_port_rf[0];
  /* vlm5030_gl.vhd:1481:73  */
  assign n14382_o = n14380_o | n14381_o;
  /* vlm5030_gl.vhd:1481:97  */
  assign n14383_o = addshift_block_cin[0];
  /* vlm5030_gl.vhd:1481:90  */
  assign n14384_o = n14382_o & n14383_o;
  /* vlm5030_gl.vhd:1481:54  */
  assign n14385_o = n14379_o | n14384_o;
  assign n14388_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14395_o = c2d4[1];
  /* vlm5030_gl.vhd:1489:31  */
  assign n14396_o = addshift_block_sum[0];
  /* vlm5030_gl.vhd:1496:27  */
  assign n14402_o = addshift_block_cin[10];
  /* vlm5030_gl.vhd:1496:52  */
  assign n14403_o = addshift_block_port_nid[9];
  /* vlm5030_gl.vhd:1496:40  */
  assign n14404_o = n14402_o ^ n14403_o;
  /* vlm5030_gl.vhd:1496:74  */
  assign n14405_o = addshift_block_port_rf[9];
  /* vlm5030_gl.vhd:1496:63  */
  assign n14406_o = n14404_o ^ n14405_o;
  assign n14409_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14416_o = c2d4[1];
  /* vlm5030_gl.vhd:1501:36  */
  assign n14417_o = addshift_block_sum[10];
  /* vlm5030_gl.vhd:1505:33  */
  assign n14423_o = addshift_block_sumlat[10];
  /* vlm5030_gl.vhd:1507:17  */
  assign n14424_o = addshift_block_sum[9:0];
  assign n14425_o = addshift_block_nidlat[0];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14426_o = n14348_o ? n14349_o : n14425_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n14341_o)
    n14427_q <= n14426_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14428_o = addshift_block_nidlat[1];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14429_o = n14285_o ? n14286_o : n14428_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n14278_o)
    n14430_q <= n14429_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14431_o = addshift_block_nidlat[2];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14432_o = n14222_o ? n14223_o : n14431_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n14215_o)
    n14433_q <= n14432_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14434_o = addshift_block_nidlat[3];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14435_o = n14159_o ? n14160_o : n14434_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n14152_o)
    n14436_q <= n14435_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14437_o = addshift_block_nidlat[4];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14438_o = n14096_o ? n14097_o : n14437_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n14089_o)
    n14439_q <= n14438_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14440_o = addshift_block_nidlat[5];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14441_o = n14033_o ? n14034_o : n14440_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n14026_o)
    n14442_q <= n14441_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14443_o = addshift_block_nidlat[6];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14444_o = n13970_o ? n13971_o : n14443_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n13963_o)
    n14445_q <= n14444_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14446_o = addshift_block_nidlat[7];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14447_o = n13907_o ? n13908_o : n14446_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n13900_o)
    n14448_q <= n14447_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14449_o = addshift_block_nidlat[8];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14450_o = n13844_o ? n13845_o : n14449_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n13837_o)
    n14451_q <= n14450_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14452_o = addshift_block_nidlat[9];
  /* vlm5030_gl.vhd:1465:9  */
  assign n14453_o = n13781_o ? n13782_o : n14452_o;
  /* vlm5030_gl.vhd:1465:9  */
  always @(posedge n13774_o)
    n14454_q <= n14453_o;
  /* vlm5030_gl.vhd:1465:9  */
  assign n14455_o = {n14454_q, n14451_q, n14448_q, n14445_q, n14442_q, n14439_q, n14436_q, n14433_q, n14430_q, n14427_q};
  assign n14456_o = {n13790_o, n13853_o, n13916_o, n13979_o, n14042_o, n14105_o, n14168_o, n14231_o, n14294_o, n14357_o};
  assign n14457_o = {n13800_o, n13863_o, n13926_o, n13989_o, n14052_o, n14115_o, n14178_o, n14241_o, n14304_o, n14367_o};
  assign n14458_o = addshift_block_sumlat[10];
  /* vlm5030_gl.vhd:1499:7  */
  assign n14459_o = n14416_o ? n14417_o : n14458_o;
  /* vlm5030_gl.vhd:1499:7  */
  always @(posedge n14409_o)
    n14460_q <= n14459_o;
  /* vlm5030_gl.vhd:1499:7  */
  assign n14461_o = addshift_block_sumlat[0];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14462_o = n14395_o ? n14396_o : n14461_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n14388_o)
    n14463_q <= n14462_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14464_o = addshift_block_sumlat[1];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14465_o = n14332_o ? n14333_o : n14464_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n14325_o)
    n14466_q <= n14465_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14467_o = addshift_block_sumlat[2];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14468_o = n14269_o ? n14270_o : n14467_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n14262_o)
    n14469_q <= n14468_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14470_o = addshift_block_sumlat[3];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14471_o = n14206_o ? n14207_o : n14470_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n14199_o)
    n14472_q <= n14471_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14473_o = addshift_block_sumlat[4];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14474_o = n14143_o ? n14144_o : n14473_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n14136_o)
    n14475_q <= n14474_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14476_o = addshift_block_sumlat[5];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14477_o = n14080_o ? n14081_o : n14476_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n14073_o)
    n14478_q <= n14477_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14479_o = addshift_block_sumlat[6];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14480_o = n14017_o ? n14018_o : n14479_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n14010_o)
    n14481_q <= n14480_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14482_o = addshift_block_sumlat[7];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14483_o = n13954_o ? n13955_o : n14482_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n13947_o)
    n14484_q <= n14483_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14485_o = addshift_block_sumlat[8];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14486_o = n13891_o ? n13892_o : n14485_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n13884_o)
    n14487_q <= n14486_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14488_o = addshift_block_sumlat[9];
  /* vlm5030_gl.vhd:1487:9  */
  assign n14489_o = n13828_o ? n13829_o : n14488_o;
  /* vlm5030_gl.vhd:1487:9  */
  always @(posedge n13821_o)
    n14490_q <= n14489_o;
  /* vlm5030_gl.vhd:1487:9  */
  assign n14491_o = {n14423_o, n14460_q, n14490_q, n14487_q, n14484_q, n14481_q, n14478_q, n14475_q, n14472_q, n14469_q, n14466_q, n14463_q};
  assign n14492_o = {n13818_o, n13881_o, n13944_o, n14007_o, n14070_o, n14133_o, n14196_o, n14259_o, n14322_o, n14385_o, n13771_o};
  assign n14493_o = {n14406_o, n13809_o, n13872_o, n13935_o, n13998_o, n14061_o, n14124_o, n14187_o, n14250_o, n14313_o, n14376_o};
  /* vlm5030_gl.vhd:1517:12  */
  always @*
    pitchinc_block_pitchlat = n14624_q; // (isignal)
  initial
    pitchinc_block_pitchlat = 7'b0000000;
  /* vlm5030_gl.vhd:1518:11  */
  always @*
    pitchinc_block_pitchreg = n14626_q; // (isignal)
  initial
    pitchinc_block_pitchreg = 7'b0000000;
  /* vlm5030_gl.vhd:1519:12  */
  assign pitchinc_block_toggle = n14627_o; // (signal)
  /* clock_functions_pack.vhd:116:26  */
  assign n14502_o = c2d4[0];
  /* clock_functions_pack.vhd:117:26  */
  assign n14503_o = c2d4[1];
  /* clock_functions_pack.vhd:117:30  */
  assign n14504_o = ~(n14503_o & updtpitch);
  /* clock_functions_pack.vhd:118:26  */
  assign n14505_o = c2d4[3];
  /* clock_functions_pack.vhd:118:31  */
  assign n14506_o = n14505_o & updtpitch;
  /* clock_functions_pack.vhd:119:26  */
  assign n14507_o = c2d4[2];
  /* clock_functions_pack.vhd:119:31  */
  assign n14508_o = n14507_o & updtpitch;
  assign n14509_o = {n14508_o, n14506_o, n14504_o, n14502_o};
  /* clock_functions_pack.vhd:75:25  */
  assign n14514_o = n14509_o[0];
  /* clock_functions_pack.vhd:76:29  */
  assign n14515_o = n14509_o[1];
  /* clock_functions_pack.vhd:76:21  */
  assign n14516_o = ~n14515_o;
  /* clock_functions_pack.vhd:77:25  */
  assign n14517_o = n14509_o[3];
  /* clock_functions_pack.vhd:78:25  */
  assign n14518_o = n14509_o[2];
  assign n14519_o = {n14518_o, n14517_o, n14516_o, n14514_o};
  assign n14522_o = osc[0];
  /* clock_functions_pack.vhd:175:17  */
  assign n14529_o = enpitchlat[1];
  /* vlm5030_gl.vhd:1528:26  */
  assign n14530_o = nid[9:3];
  assign n14541_o = clk2ena[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n14543_o = clk2ena[2];
  /* vlm5030_gl.vhd:1545:22  */
  assign n14545_o = pitchinc_block_toggle[6];
  /* vlm5030_gl.vhd:1546:44  */
  assign n14546_o = pitchinc_block_pitchreg[6];
  /* vlm5030_gl.vhd:1546:32  */
  assign n14547_o = ~n14546_o;
  assign n14548_o = pitchinc_block_pitchreg[6];
  /* vlm5030_gl.vhd:1545:13  */
  assign n14549_o = n14545_o ? n14547_o : n14548_o;
  /* vlm5030_gl.vhd:1545:22  */
  assign n14550_o = pitchinc_block_toggle[5];
  /* vlm5030_gl.vhd:1546:44  */
  assign n14551_o = pitchinc_block_pitchreg[5];
  /* vlm5030_gl.vhd:1546:32  */
  assign n14552_o = ~n14551_o;
  assign n14553_o = pitchinc_block_pitchreg[5];
  /* vlm5030_gl.vhd:1545:13  */
  assign n14554_o = n14550_o ? n14552_o : n14553_o;
  /* vlm5030_gl.vhd:1545:22  */
  assign n14555_o = pitchinc_block_toggle[4];
  /* vlm5030_gl.vhd:1546:44  */
  assign n14556_o = pitchinc_block_pitchreg[4];
  /* vlm5030_gl.vhd:1546:32  */
  assign n14557_o = ~n14556_o;
  assign n14558_o = pitchinc_block_pitchreg[4];
  /* vlm5030_gl.vhd:1545:13  */
  assign n14559_o = n14555_o ? n14557_o : n14558_o;
  /* vlm5030_gl.vhd:1545:22  */
  assign n14560_o = pitchinc_block_toggle[3];
  /* vlm5030_gl.vhd:1546:44  */
  assign n14561_o = pitchinc_block_pitchreg[3];
  /* vlm5030_gl.vhd:1546:32  */
  assign n14562_o = ~n14561_o;
  assign n14563_o = pitchinc_block_pitchreg[3];
  /* vlm5030_gl.vhd:1545:13  */
  assign n14564_o = n14560_o ? n14562_o : n14563_o;
  /* vlm5030_gl.vhd:1545:22  */
  assign n14565_o = pitchinc_block_toggle[2];
  /* vlm5030_gl.vhd:1546:44  */
  assign n14566_o = pitchinc_block_pitchreg[2];
  /* vlm5030_gl.vhd:1546:32  */
  assign n14567_o = ~n14566_o;
  assign n14568_o = pitchinc_block_pitchreg[2];
  /* vlm5030_gl.vhd:1545:13  */
  assign n14569_o = n14565_o ? n14567_o : n14568_o;
  /* vlm5030_gl.vhd:1545:22  */
  assign n14570_o = pitchinc_block_toggle[1];
  /* vlm5030_gl.vhd:1546:44  */
  assign n14571_o = pitchinc_block_pitchreg[1];
  /* vlm5030_gl.vhd:1546:32  */
  assign n14572_o = ~n14571_o;
  assign n14573_o = pitchinc_block_pitchreg[1];
  /* vlm5030_gl.vhd:1545:13  */
  assign n14574_o = n14570_o ? n14572_o : n14573_o;
  /* vlm5030_gl.vhd:1545:22  */
  assign n14575_o = pitchinc_block_toggle[0];
  /* vlm5030_gl.vhd:1546:44  */
  assign n14576_o = pitchinc_block_pitchreg[0];
  /* vlm5030_gl.vhd:1546:32  */
  assign n14577_o = ~n14576_o;
  assign n14578_o = pitchinc_block_pitchreg[0];
  /* vlm5030_gl.vhd:1545:13  */
  assign n14579_o = n14575_o ? n14577_o : n14578_o;
  assign n14580_o = {n14549_o, n14554_o, n14559_o, n14564_o, n14569_o, n14574_o, n14579_o};
  /* vlm5030_gl.vhd:1539:9  */
  assign n14581_o = pitchoverflow ? pitchinc_block_pitchlat : n14580_o;
  /* vlm5030_gl.vhd:1556:35  */
  assign n14587_o = pitchinc_block_pitchreg[0];
  /* vlm5030_gl.vhd:1556:23  */
  assign n14588_o = ~n14587_o;
  /* vlm5030_gl.vhd:1556:59  */
  assign n14589_o = pitchinc_block_toggle[0];
  /* vlm5030_gl.vhd:1556:49  */
  assign n14590_o = ~n14589_o;
  /* vlm5030_gl.vhd:1556:44  */
  assign n14591_o = ~(n14588_o | n14590_o);
  /* vlm5030_gl.vhd:1556:35  */
  assign n14592_o = pitchinc_block_pitchreg[1];
  /* vlm5030_gl.vhd:1556:23  */
  assign n14593_o = ~n14592_o;
  /* vlm5030_gl.vhd:1556:59  */
  assign n14594_o = pitchinc_block_toggle[1];
  /* vlm5030_gl.vhd:1556:49  */
  assign n14595_o = ~n14594_o;
  /* vlm5030_gl.vhd:1556:44  */
  assign n14596_o = ~(n14593_o | n14595_o);
  /* vlm5030_gl.vhd:1556:35  */
  assign n14597_o = pitchinc_block_pitchreg[2];
  /* vlm5030_gl.vhd:1556:23  */
  assign n14598_o = ~n14597_o;
  /* vlm5030_gl.vhd:1556:59  */
  assign n14599_o = pitchinc_block_toggle[2];
  /* vlm5030_gl.vhd:1556:49  */
  assign n14600_o = ~n14599_o;
  /* vlm5030_gl.vhd:1556:44  */
  assign n14601_o = ~(n14598_o | n14600_o);
  /* vlm5030_gl.vhd:1556:35  */
  assign n14602_o = pitchinc_block_pitchreg[3];
  /* vlm5030_gl.vhd:1556:23  */
  assign n14603_o = ~n14602_o;
  /* vlm5030_gl.vhd:1556:59  */
  assign n14604_o = pitchinc_block_toggle[3];
  /* vlm5030_gl.vhd:1556:49  */
  assign n14605_o = ~n14604_o;
  /* vlm5030_gl.vhd:1556:44  */
  assign n14606_o = ~(n14603_o | n14605_o);
  /* vlm5030_gl.vhd:1556:35  */
  assign n14607_o = pitchinc_block_pitchreg[4];
  /* vlm5030_gl.vhd:1556:23  */
  assign n14608_o = ~n14607_o;
  /* vlm5030_gl.vhd:1556:59  */
  assign n14609_o = pitchinc_block_toggle[4];
  /* vlm5030_gl.vhd:1556:49  */
  assign n14610_o = ~n14609_o;
  /* vlm5030_gl.vhd:1556:44  */
  assign n14611_o = ~(n14608_o | n14610_o);
  /* vlm5030_gl.vhd:1556:35  */
  assign n14612_o = pitchinc_block_pitchreg[5];
  /* vlm5030_gl.vhd:1556:23  */
  assign n14613_o = ~n14612_o;
  /* vlm5030_gl.vhd:1556:59  */
  assign n14614_o = pitchinc_block_toggle[5];
  /* vlm5030_gl.vhd:1556:49  */
  assign n14615_o = ~n14614_o;
  /* vlm5030_gl.vhd:1556:44  */
  assign n14616_o = ~(n14613_o | n14615_o);
  /* vlm5030_gl.vhd:1556:35  */
  assign n14617_o = pitchinc_block_pitchreg[6];
  /* vlm5030_gl.vhd:1556:23  */
  assign n14618_o = ~n14617_o;
  /* vlm5030_gl.vhd:1556:59  */
  assign n14619_o = pitchinc_block_toggle[6];
  /* vlm5030_gl.vhd:1556:49  */
  assign n14620_o = ~n14619_o;
  /* vlm5030_gl.vhd:1556:44  */
  assign n14621_o = ~(n14618_o | n14620_o);
  /* vlm5030_gl.vhd:1559:28  */
  assign n14622_o = pitchinc_block_toggle[7];
  /* vlm5030_gl.vhd:1526:7  */
  assign n14623_o = n14529_o ? n14530_o : pitchinc_block_pitchlat;
  /* vlm5030_gl.vhd:1526:7  */
  always @(posedge n14522_o)
    n14624_q <= n14623_o;
  initial
    n14624_q = 7'b0000000;
  /* vlm5030_gl.vhd:1538:7  */
  assign n14625_o = n14543_o ? n14581_o : pitchinc_block_pitchreg;
  /* vlm5030_gl.vhd:1538:7  */
  always @(posedge n14541_o or posedge rstdel)
    if (rstdel)
      n14626_q <= 7'b0000000;
    else
      n14626_q <= n14625_o;
  /* vlm5030_gl.vhd:1535:7  */
  assign n14627_o = {n14621_o, n14616_o, n14611_o, n14606_o, n14601_o, n14596_o, n14591_o, 1'b1};
  /* vlm5030_gl.vhd:1564:27  */
  assign n14629_o = dq[6];
  /* vlm5030_gl.vhd:1564:37  */
  assign n14630_o = dq[7];
  /* vlm5030_gl.vhd:1564:31  */
  assign n14631_o = n14629_o ^ n14630_o;
  /* vlm5030_gl.vhd:1564:21  */
  assign n14632_o = ~n14631_o;
  /* vlm5030_gl.vhd:1564:43  */
  assign n14633_o = n14632_o | tstend2id;
  /* clock_functions_pack.vhd:147:24  */
  assign n14638_o = nc2d1[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n14639_o = n14633_o | n14638_o;
  /* vlm5030_gl.vhd:1564:15  */
  assign n14640_o = ~n14639_o;
  /* vlm5030_gl.vhd:1572:12  */
  assign nid_block_wl = n14645_o; // (signal)
  /* vlm5030_gl.vhd:1575:34  */
  assign n14641_o = {tstend2id, enrf2id};
  /* vlm5030_gl.vhd:1575:44  */
  assign n14642_o = {n14641_o, ensum2id};
  /* vlm5030_gl.vhd:1575:55  */
  assign n14643_o = {n14642_o, updtpitch};
  /* vlm5030_gl.vhd:1575:67  */
  assign n14644_o = {n14643_o, enidlinv2id};
  /* vlm5030_gl.vhd:1575:82  */
  assign n14645_o = {n14644_o, enmem02id};
  /* vlm5030_gl.vhd:1577:28  */
  assign n14647_o = i_d[0];
  /* vlm5030_gl.vhd:1577:40  */
  assign n14648_o = rfdo[0];
  /* vlm5030_gl.vhd:1577:34  */
  assign n14649_o = {n14647_o, n14648_o};
  /* vlm5030_gl.vhd:1577:51  */
  assign n14650_o = assum[0];
  /* vlm5030_gl.vhd:1577:44  */
  assign n14651_o = {n14649_o, n14650_o};
  /* vlm5030_gl.vhd:1577:55  */
  assign n14653_o = {n14651_o, 1'b0};
  /* vlm5030_gl.vhd:1577:78  */
  assign n14654_o = idlat[0];
  /* vlm5030_gl.vhd:1577:69  */
  assign n14655_o = ~n14654_o;
  /* vlm5030_gl.vhd:1577:67  */
  assign n14656_o = {n14653_o, n14655_o};
  /* vlm5030_gl.vhd:1577:91  */
  assign n14657_o = nmem0do[0];
  /* vlm5030_gl.vhd:1577:82  */
  assign n14658_o = {n14656_o, n14657_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n14664_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n14665_o = n14658_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n14666_o = n14664_o & n14665_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14668_o = 1'b0 | n14666_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14670_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n14671_o = n14658_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n14672_o = n14670_o & n14671_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14673_o = n14668_o | n14672_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14674_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n14675_o = n14658_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n14676_o = n14674_o & n14675_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14677_o = n14673_o | n14676_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14678_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n14679_o = n14658_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n14680_o = n14678_o & n14679_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14681_o = n14677_o | n14680_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14682_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n14683_o = n14658_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n14684_o = n14682_o & n14683_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14685_o = n14681_o | n14684_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14686_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n14687_o = n14658_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n14688_o = n14686_o & n14687_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14689_o = n14685_o | n14688_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n14690_o = ~n14689_o;
  /* vlm5030_gl.vhd:1578:28  */
  assign n14692_o = i_d[1];
  /* vlm5030_gl.vhd:1578:40  */
  assign n14693_o = rfdo[1];
  /* vlm5030_gl.vhd:1578:34  */
  assign n14694_o = {n14692_o, n14693_o};
  /* vlm5030_gl.vhd:1578:51  */
  assign n14695_o = assum[1];
  /* vlm5030_gl.vhd:1578:44  */
  assign n14696_o = {n14694_o, n14695_o};
  /* vlm5030_gl.vhd:1578:55  */
  assign n14698_o = {n14696_o, 1'b0};
  /* vlm5030_gl.vhd:1578:78  */
  assign n14699_o = idlat[1];
  /* vlm5030_gl.vhd:1578:69  */
  assign n14700_o = ~n14699_o;
  /* vlm5030_gl.vhd:1578:67  */
  assign n14701_o = {n14698_o, n14700_o};
  /* vlm5030_gl.vhd:1578:91  */
  assign n14702_o = nmem0do[1];
  /* vlm5030_gl.vhd:1578:82  */
  assign n14703_o = {n14701_o, n14702_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n14709_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n14710_o = n14703_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n14711_o = n14709_o & n14710_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14713_o = 1'b0 | n14711_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14715_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n14716_o = n14703_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n14717_o = n14715_o & n14716_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14718_o = n14713_o | n14717_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14719_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n14720_o = n14703_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n14721_o = n14719_o & n14720_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14722_o = n14718_o | n14721_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14723_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n14724_o = n14703_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n14725_o = n14723_o & n14724_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14726_o = n14722_o | n14725_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14727_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n14728_o = n14703_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n14729_o = n14727_o & n14728_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14730_o = n14726_o | n14729_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14731_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n14732_o = n14703_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n14733_o = n14731_o & n14732_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14734_o = n14730_o | n14733_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n14735_o = ~n14734_o;
  /* vlm5030_gl.vhd:1579:28  */
  assign n14737_o = i_d[2];
  /* vlm5030_gl.vhd:1579:40  */
  assign n14738_o = rfdo[2];
  /* vlm5030_gl.vhd:1579:34  */
  assign n14739_o = {n14737_o, n14738_o};
  /* vlm5030_gl.vhd:1579:51  */
  assign n14740_o = assum[2];
  /* vlm5030_gl.vhd:1579:44  */
  assign n14741_o = {n14739_o, n14740_o};
  /* vlm5030_gl.vhd:1579:55  */
  assign n14743_o = {n14741_o, 1'b0};
  /* vlm5030_gl.vhd:1579:78  */
  assign n14744_o = idlat[2];
  /* vlm5030_gl.vhd:1579:69  */
  assign n14745_o = ~n14744_o;
  /* vlm5030_gl.vhd:1579:67  */
  assign n14746_o = {n14743_o, n14745_o};
  /* vlm5030_gl.vhd:1579:91  */
  assign n14747_o = nmem0do[2];
  /* vlm5030_gl.vhd:1579:82  */
  assign n14748_o = {n14746_o, n14747_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n14754_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n14755_o = n14748_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n14756_o = n14754_o & n14755_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14758_o = 1'b0 | n14756_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14760_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n14761_o = n14748_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n14762_o = n14760_o & n14761_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14763_o = n14758_o | n14762_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14764_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n14765_o = n14748_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n14766_o = n14764_o & n14765_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14767_o = n14763_o | n14766_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14768_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n14769_o = n14748_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n14770_o = n14768_o & n14769_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14771_o = n14767_o | n14770_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14772_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n14773_o = n14748_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n14774_o = n14772_o & n14773_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14775_o = n14771_o | n14774_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14776_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n14777_o = n14748_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n14778_o = n14776_o & n14777_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14779_o = n14775_o | n14778_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n14780_o = ~n14779_o;
  /* vlm5030_gl.vhd:1580:28  */
  assign n14782_o = i_d[3];
  /* vlm5030_gl.vhd:1580:40  */
  assign n14783_o = rfdo[3];
  /* vlm5030_gl.vhd:1580:34  */
  assign n14784_o = {n14782_o, n14783_o};
  /* vlm5030_gl.vhd:1580:51  */
  assign n14785_o = assum[3];
  /* vlm5030_gl.vhd:1580:44  */
  assign n14786_o = {n14784_o, n14785_o};
  /* vlm5030_gl.vhd:1580:55  */
  assign n14788_o = {n14786_o, 1'b0};
  /* vlm5030_gl.vhd:1580:78  */
  assign n14789_o = idlat[3];
  /* vlm5030_gl.vhd:1580:69  */
  assign n14790_o = ~n14789_o;
  /* vlm5030_gl.vhd:1580:67  */
  assign n14791_o = {n14788_o, n14790_o};
  /* vlm5030_gl.vhd:1580:91  */
  assign n14792_o = nmem0do[3];
  /* vlm5030_gl.vhd:1580:82  */
  assign n14793_o = {n14791_o, n14792_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n14799_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n14800_o = n14793_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n14801_o = n14799_o & n14800_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14803_o = 1'b0 | n14801_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14805_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n14806_o = n14793_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n14807_o = n14805_o & n14806_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14808_o = n14803_o | n14807_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14809_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n14810_o = n14793_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n14811_o = n14809_o & n14810_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14812_o = n14808_o | n14811_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14813_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n14814_o = n14793_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n14815_o = n14813_o & n14814_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14816_o = n14812_o | n14815_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14817_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n14818_o = n14793_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n14819_o = n14817_o & n14818_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14820_o = n14816_o | n14819_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14821_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n14822_o = n14793_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n14823_o = n14821_o & n14822_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14824_o = n14820_o | n14823_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n14825_o = ~n14824_o;
  /* vlm5030_gl.vhd:1581:28  */
  assign n14827_o = i_d[4];
  /* vlm5030_gl.vhd:1581:40  */
  assign n14828_o = rfdo[4];
  /* vlm5030_gl.vhd:1581:34  */
  assign n14829_o = {n14827_o, n14828_o};
  /* vlm5030_gl.vhd:1581:51  */
  assign n14830_o = assum[4];
  /* vlm5030_gl.vhd:1581:44  */
  assign n14831_o = {n14829_o, n14830_o};
  /* vlm5030_gl.vhd:1581:55  */
  assign n14833_o = {n14831_o, 1'b0};
  /* vlm5030_gl.vhd:1581:78  */
  assign n14834_o = idlat[4];
  /* vlm5030_gl.vhd:1581:69  */
  assign n14835_o = ~n14834_o;
  /* vlm5030_gl.vhd:1581:67  */
  assign n14836_o = {n14833_o, n14835_o};
  /* vlm5030_gl.vhd:1581:91  */
  assign n14837_o = nmem0do[4];
  /* vlm5030_gl.vhd:1581:82  */
  assign n14838_o = {n14836_o, n14837_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n14844_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n14845_o = n14838_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n14846_o = n14844_o & n14845_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14848_o = 1'b0 | n14846_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14850_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n14851_o = n14838_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n14852_o = n14850_o & n14851_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14853_o = n14848_o | n14852_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14854_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n14855_o = n14838_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n14856_o = n14854_o & n14855_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14857_o = n14853_o | n14856_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14858_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n14859_o = n14838_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n14860_o = n14858_o & n14859_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14861_o = n14857_o | n14860_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14862_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n14863_o = n14838_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n14864_o = n14862_o & n14863_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14865_o = n14861_o | n14864_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14866_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n14867_o = n14838_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n14868_o = n14866_o & n14867_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14869_o = n14865_o | n14868_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n14870_o = ~n14869_o;
  /* vlm5030_gl.vhd:1582:28  */
  assign n14872_o = i_d[5];
  /* vlm5030_gl.vhd:1582:40  */
  assign n14873_o = rfdo[5];
  /* vlm5030_gl.vhd:1582:34  */
  assign n14874_o = {n14872_o, n14873_o};
  /* vlm5030_gl.vhd:1582:51  */
  assign n14875_o = assum[5];
  /* vlm5030_gl.vhd:1582:44  */
  assign n14876_o = {n14874_o, n14875_o};
  /* vlm5030_gl.vhd:1582:55  */
  assign n14878_o = {n14876_o, 1'b0};
  /* vlm5030_gl.vhd:1582:78  */
  assign n14879_o = idlat[5];
  /* vlm5030_gl.vhd:1582:69  */
  assign n14880_o = ~n14879_o;
  /* vlm5030_gl.vhd:1582:67  */
  assign n14881_o = {n14878_o, n14880_o};
  /* vlm5030_gl.vhd:1582:91  */
  assign n14882_o = nmem0do[5];
  /* vlm5030_gl.vhd:1582:82  */
  assign n14883_o = {n14881_o, n14882_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n14889_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n14890_o = n14883_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n14891_o = n14889_o & n14890_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14893_o = 1'b0 | n14891_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14895_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n14896_o = n14883_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n14897_o = n14895_o & n14896_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14898_o = n14893_o | n14897_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14899_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n14900_o = n14883_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n14901_o = n14899_o & n14900_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14902_o = n14898_o | n14901_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14903_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n14904_o = n14883_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n14905_o = n14903_o & n14904_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14906_o = n14902_o | n14905_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14907_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n14908_o = n14883_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n14909_o = n14907_o & n14908_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14910_o = n14906_o | n14909_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14911_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n14912_o = n14883_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n14913_o = n14911_o & n14912_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14914_o = n14910_o | n14913_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n14915_o = ~n14914_o;
  /* vlm5030_gl.vhd:1583:28  */
  assign n14917_o = i_d[6];
  /* vlm5030_gl.vhd:1583:40  */
  assign n14918_o = rfdo[6];
  /* vlm5030_gl.vhd:1583:34  */
  assign n14919_o = {n14917_o, n14918_o};
  /* vlm5030_gl.vhd:1583:51  */
  assign n14920_o = assum[6];
  /* vlm5030_gl.vhd:1583:44  */
  assign n14921_o = {n14919_o, n14920_o};
  /* vlm5030_gl.vhd:1583:55  */
  assign n14922_o = {n14921_o, pitchmod};
  /* vlm5030_gl.vhd:1583:78  */
  assign n14923_o = idlat[6];
  /* vlm5030_gl.vhd:1583:69  */
  assign n14924_o = ~n14923_o;
  /* vlm5030_gl.vhd:1583:67  */
  assign n14925_o = {n14922_o, n14924_o};
  /* vlm5030_gl.vhd:1583:91  */
  assign n14926_o = nmem0do[6];
  /* vlm5030_gl.vhd:1583:82  */
  assign n14927_o = {n14925_o, n14926_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n14933_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n14934_o = n14927_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n14935_o = n14933_o & n14934_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14937_o = 1'b0 | n14935_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14939_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n14940_o = n14927_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n14941_o = n14939_o & n14940_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14942_o = n14937_o | n14941_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14943_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n14944_o = n14927_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n14945_o = n14943_o & n14944_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14946_o = n14942_o | n14945_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14947_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n14948_o = n14927_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n14949_o = n14947_o & n14948_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14950_o = n14946_o | n14949_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14951_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n14952_o = n14927_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n14953_o = n14951_o & n14952_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14954_o = n14950_o | n14953_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14955_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n14956_o = n14927_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n14957_o = n14955_o & n14956_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14958_o = n14954_o | n14957_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n14959_o = ~n14958_o;
  /* vlm5030_gl.vhd:1584:28  */
  assign n14961_o = i_d[7];
  /* vlm5030_gl.vhd:1584:40  */
  assign n14962_o = rfdo[7];
  /* vlm5030_gl.vhd:1584:34  */
  assign n14963_o = {n14961_o, n14962_o};
  /* vlm5030_gl.vhd:1584:51  */
  assign n14964_o = assum[7];
  /* vlm5030_gl.vhd:1584:44  */
  assign n14965_o = {n14963_o, n14964_o};
  /* vlm5030_gl.vhd:1584:55  */
  assign n14967_o = {n14965_o, 1'b0};
  /* vlm5030_gl.vhd:1584:78  */
  assign n14968_o = idlat[7];
  /* vlm5030_gl.vhd:1584:69  */
  assign n14969_o = ~n14968_o;
  /* vlm5030_gl.vhd:1584:67  */
  assign n14970_o = {n14967_o, n14969_o};
  /* vlm5030_gl.vhd:1584:91  */
  assign n14971_o = nmem0do[7];
  /* vlm5030_gl.vhd:1584:82  */
  assign n14972_o = {n14970_o, n14971_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n14978_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n14979_o = n14972_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n14980_o = n14978_o & n14979_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14982_o = 1'b0 | n14980_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14984_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n14985_o = n14972_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n14986_o = n14984_o & n14985_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14987_o = n14982_o | n14986_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14988_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n14989_o = n14972_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n14990_o = n14988_o & n14989_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14991_o = n14987_o | n14990_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14992_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n14993_o = n14972_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n14994_o = n14992_o & n14993_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14995_o = n14991_o | n14994_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n14996_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n14997_o = n14972_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n14998_o = n14996_o & n14997_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n14999_o = n14995_o | n14998_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15000_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15001_o = n14972_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15002_o = n15000_o & n15001_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15003_o = n14999_o | n15002_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15004_o = ~n15003_o;
  /* vlm5030_gl.vhd:1585:28  */
  assign n15006_o = i_d[0];
  /* vlm5030_gl.vhd:1585:40  */
  assign n15007_o = rfdo[8];
  /* vlm5030_gl.vhd:1585:34  */
  assign n15008_o = {n15006_o, n15007_o};
  /* vlm5030_gl.vhd:1585:51  */
  assign n15009_o = assum[8];
  /* vlm5030_gl.vhd:1585:44  */
  assign n15010_o = {n15008_o, n15009_o};
  /* vlm5030_gl.vhd:1585:55  */
  assign n15012_o = {n15010_o, 1'b0};
  /* vlm5030_gl.vhd:1585:67  */
  assign n15014_o = {n15012_o, 1'b0};
  /* vlm5030_gl.vhd:1585:91  */
  assign n15015_o = nmem0do[8];
  /* vlm5030_gl.vhd:1585:82  */
  assign n15016_o = {n15014_o, n15015_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15022_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n15023_o = n15016_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n15024_o = n15022_o & n15023_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15026_o = 1'b0 | n15024_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15028_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n15029_o = n15016_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n15030_o = n15028_o & n15029_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15031_o = n15026_o | n15030_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15032_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n15033_o = n15016_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n15034_o = n15032_o & n15033_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15035_o = n15031_o | n15034_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15036_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n15037_o = n15016_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n15038_o = n15036_o & n15037_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15039_o = n15035_o | n15038_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15040_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15041_o = n15016_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15042_o = n15040_o & n15041_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15043_o = n15039_o | n15042_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15044_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15045_o = n15016_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15046_o = n15044_o & n15045_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15047_o = n15043_o | n15046_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15048_o = ~n15047_o;
  /* vlm5030_gl.vhd:1586:28  */
  assign n15050_o = i_d[1];
  /* vlm5030_gl.vhd:1586:40  */
  assign n15051_o = rfdo[9];
  /* vlm5030_gl.vhd:1586:34  */
  assign n15052_o = {n15050_o, n15051_o};
  /* vlm5030_gl.vhd:1586:51  */
  assign n15053_o = assum[9];
  /* vlm5030_gl.vhd:1586:44  */
  assign n15054_o = {n15052_o, n15053_o};
  /* vlm5030_gl.vhd:1586:55  */
  assign n15056_o = {n15054_o, 1'b0};
  /* vlm5030_gl.vhd:1586:67  */
  assign n15058_o = {n15056_o, 1'b0};
  /* vlm5030_gl.vhd:1586:91  */
  assign n15059_o = nmem0do[9];
  /* vlm5030_gl.vhd:1586:82  */
  assign n15060_o = {n15058_o, n15059_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15066_o = nid_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n15067_o = n15060_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n15068_o = n15066_o & n15067_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15070_o = 1'b0 | n15068_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15072_o = nid_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n15073_o = n15060_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n15074_o = n15072_o & n15073_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15075_o = n15070_o | n15074_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15076_o = nid_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n15077_o = n15060_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n15078_o = n15076_o & n15077_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15079_o = n15075_o | n15078_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15080_o = nid_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n15081_o = n15060_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n15082_o = n15080_o & n15081_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15083_o = n15079_o | n15082_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15084_o = nid_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15085_o = n15060_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15086_o = n15084_o & n15085_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15087_o = n15083_o | n15086_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15088_o = nid_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15089_o = n15060_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15090_o = n15088_o & n15089_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15091_o = n15087_o | n15090_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15092_o = ~n15091_o;
  /* vlm5030_gl.vhd:1596:12  */
  assign idlat_block_idlaten = n15105_o; // (signal)
  /* vlm5030_gl.vhd:1597:12  */
  assign idlat_block_n = n15124_o; // (signal)
  /* vlm5030_gl.vhd:1600:37  */
  assign n15094_o = fsromdo[6];
  /* vlm5030_gl.vhd:1600:26  */
  assign n15095_o = ~n15094_o;
  /* vlm5030_gl.vhd:1600:56  */
  assign n15096_o = xromdo[10];
  /* vlm5030_gl.vhd:1600:46  */
  assign n15097_o = ~n15096_o;
  /* vlm5030_gl.vhd:1600:42  */
  assign n15098_o = n15095_o | n15097_o;
  /* clock_functions_pack.vhd:147:24  */
  assign n15103_o = nc2d8[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n15104_o = n15098_o | n15103_o;
  /* vlm5030_gl.vhd:1600:20  */
  assign n15105_o = ~n15104_o;
  /* vlm5030_gl.vhd:1601:36  */
  assign n15107_o = xromdo[10];
  /* vlm5030_gl.vhd:1601:26  */
  assign n15108_o = ~n15107_o;
  /* vlm5030_gl.vhd:1601:42  */
  assign n15109_o = n15108_o | tstend2id;
  /* clock_functions_pack.vhd:147:24  */
  assign n15114_o = nc2d1[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n15115_o = n15109_o | n15114_o;
  /* vlm5030_gl.vhd:1601:20  */
  assign n15116_o = ~n15115_o;
  /* vlm5030_gl.vhd:1603:29  */
  assign n15118_o = xromdo7q | tstend2ie;
  /* clock_functions_pack.vhd:147:24  */
  assign n15123_o = c2d7fin[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n15124_o = n15118_o | n15123_o;
  /* vlm5030_gl.vhd:1604:36  */
  assign n15125_o = maskdq53 & random;
  /* vlm5030_gl.vhd:1604:53  */
  assign n15126_o = ~maskdq53;
  /* vlm5030_gl.vhd:1604:67  */
  assign n15127_o = n15126_o & pitchoverflow;
  /* vlm5030_gl.vhd:1604:48  */
  assign n15128_o = n15125_o | n15127_o;
  /* vlm5030_gl.vhd:1604:21  */
  assign n15129_o = ~n15128_o;
  /* vlm5030_gl.vhd:1604:89  */
  assign n15130_o = ~(n15129_o | idlat_block_n);
  /* vlm5030_gl.vhd:1605:27  */
  assign n15131_o = idlat_block_n | random;
  /* vlm5030_gl.vhd:1605:37  */
  assign n15132_o = n15131_o | idlatall1;
  /* vlm5030_gl.vhd:1605:54  */
  assign n15133_o = ~maskdq53;
  /* vlm5030_gl.vhd:1605:50  */
  assign n15134_o = n15132_o | n15133_o;
  /* vlm5030_gl.vhd:1605:20  */
  assign n15135_o = ~n15134_o;
  assign n15138_o = osc[0];
  /* vlm5030_gl.vhd:1611:23  */
  assign n15140_o = nid[7:0];
  /* vlm5030_gl.vhd:1616:23  */
  assign n15145_o = ~idlat;
  /* vlm5030_pack.vhd:40:24  */
  assign n15151_o = n15145_o[7];
  /* vlm5030_pack.vhd:40:20  */
  assign n15153_o = 1'b0 | n15151_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n15155_o = n15145_o[6];
  /* vlm5030_pack.vhd:40:20  */
  assign n15156_o = n15153_o | n15155_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n15157_o = n15145_o[5];
  /* vlm5030_pack.vhd:40:20  */
  assign n15158_o = n15156_o | n15157_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n15159_o = n15145_o[4];
  /* vlm5030_pack.vhd:40:20  */
  assign n15160_o = n15158_o | n15159_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n15161_o = n15145_o[3];
  /* vlm5030_pack.vhd:40:20  */
  assign n15162_o = n15160_o | n15161_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n15163_o = n15145_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n15164_o = n15162_o | n15163_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n15165_o = n15145_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n15166_o = n15164_o | n15165_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n15167_o = n15145_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n15168_o = n15166_o | n15167_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n15169_o = ~n15168_o;
  /* vlm5030_gl.vhd:1626:12  */
  assign mem_block_swapa = n15320_o; // (signal)
  /* vlm5030_gl.vhd:1627:12  */
  assign mem_block_a = n15177_o; // (signal)
  /* vlm5030_gl.vhd:1629:12  */
  assign mem_block_clkmem0 = n15192_o; // (signal)
  /* vlm5030_gl.vhd:1629:21  */
  assign mem_block_clkmem1 = n15238_o; // (signal)
  /* vlm5030_gl.vhd:1629:30  */
  assign mem_block_clkmem2 = n15282_o; // (signal)
  /* vlm5030_gl.vhd:1640:27  */
  assign n15173_o = yromdo[0];
  /* vlm5030_gl.vhd:1640:27  */
  assign n15174_o = yromdo[1];
  /* vlm5030_gl.vhd:1640:27  */
  assign n15175_o = yromdo[2];
  /* vlm5030_gl.vhd:1640:27  */
  assign n15176_o = yromdo[3];
  /* vlm5030_gl.vhd:1642:10  */
  assign n15177_o = {27'b0, mem_block_swapa};  //  uext
  /* vlm5030_gl.vhd:1647:29  */
  assign n15179_o = xromdo[7];
  /* vlm5030_gl.vhd:1647:48  */
  assign n15180_o = fsromdo[6];
  /* vlm5030_gl.vhd:1647:37  */
  assign n15181_o = ~n15180_o;
  /* vlm5030_gl.vhd:1647:33  */
  assign n15182_o = n15179_o | n15181_o;
  /* vlm5030_gl.vhd:1647:76  */
  assign n15183_o = yromdo[4];
  /* vlm5030_gl.vhd:1647:66  */
  assign n15184_o = xromdo7q & n15183_o;
  /* vlm5030_gl.vhd:1647:53  */
  assign n15185_o = n15182_o | n15184_o;
  /* clock_functions_pack.vhd:147:24  */
  assign n15190_o = nc2d8[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n15191_o = n15185_o | n15190_o;
  /* vlm5030_gl.vhd:1647:18  */
  assign n15192_o = ~n15191_o;
  /* vlm5030_gl.vhd:1648:56  */
  assign n15194_o = yromdo[4];
  /* vlm5030_gl.vhd:1648:46  */
  assign n15195_o = xromdo7q & n15194_o;
  /* vlm5030_gl.vhd:1648:33  */
  assign n15196_o = tstend2id | n15195_o;
  /* clock_functions_pack.vhd:147:24  */
  assign n15201_o = nc2d1[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n15202_o = n15196_o | n15201_o;
  /* vlm5030_gl.vhd:1648:18  */
  assign n15203_o = ~n15202_o;
  assign n15205_o = osc[0];
  /* vlm5030_gl.vhd:1654:16  */
  assign n15207_o = {1'b0, mem_block_a};  //  uext
  /* vlm5030_gl.vhd:1654:16  */
  assign n15209_o = $signed(n15207_o) <= $signed(32'b00000000000000000000000000001001);
  /* vlm5030_gl.vhd:1655:18  */
  assign n15210_o = mem_block_a[3:0];  // trunc
  /* vlm5030_gl.vhd:1653:9  */
  assign n15216_o = mem_block_clkmem0 & n15209_o;
  /* vlm5030_gl.vhd:1662:25  */
  assign n15219_o = mem_block_a[3:0];  // trunc
  /* vlm5030_gl.vhd:1662:16  */
  assign n15224_o = ~n20400_data;
  /* vlm5030_gl.vhd:1662:35  */
  assign n15225_o = {1'b0, mem_block_a};  //  uext
  /* vlm5030_gl.vhd:1662:35  */
  assign n15227_o = $signed(n15225_o) <= $signed(32'b00000000000000000000000000001001);
  /* vlm5030_gl.vhd:1662:28  */
  assign n15228_o = n15227_o ? n15224_o : 10'b1111111111;
  /* vlm5030_gl.vhd:1663:16  */
  assign n15230_o = ~nmem0do;
  /* vlm5030_gl.vhd:1669:24  */
  assign n15232_o = yromdo[4];
  /* clock_functions_pack.vhd:170:25  */
  assign n15237_o = nc2d10[1];
  /* clock_functions_pack.vhd:170:16  */
  assign n15238_o = ~(n15232_o | n15237_o);
  /* vlm5030_gl.vhd:1670:29  */
  assign n15240_o = yromdo[4];
  /* vlm5030_gl.vhd:1670:33  */
  assign n15241_o = n15240_o | tstend2ie;
  /* clock_functions_pack.vhd:147:24  */
  assign n15246_o = c2d7fin[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n15247_o = n15241_o | n15246_o;
  /* vlm5030_gl.vhd:1670:18  */
  assign n15248_o = ~n15247_o;
  assign n15250_o = osc[0];
  /* vlm5030_gl.vhd:1676:16  */
  assign n15252_o = {1'b0, mem_block_a};  //  uext
  /* vlm5030_gl.vhd:1676:16  */
  assign n15254_o = $signed(n15252_o) <= $signed(32'b00000000000000000000000000001001);
  /* vlm5030_gl.vhd:1677:18  */
  assign n15255_o = mem_block_a[3:0];  // trunc
  /* vlm5030_gl.vhd:1675:9  */
  assign n15261_o = mem_block_clkmem1 & n15254_o;
  /* vlm5030_gl.vhd:1684:27  */
  assign n15264_o = mem_block_a[3:0];  // trunc
  /* vlm5030_gl.vhd:1684:18  */
  assign n15269_o = ~n20403_data;
  /* vlm5030_gl.vhd:1684:37  */
  assign n15270_o = {1'b0, mem_block_a};  //  uext
  /* vlm5030_gl.vhd:1684:37  */
  assign n15272_o = $signed(n15270_o) <= $signed(32'b00000000000000000000000000001001);
  /* vlm5030_gl.vhd:1684:30  */
  assign n15273_o = n15272_o ? n15269_o : 12'b111111111111;
  /* vlm5030_gl.vhd:1690:24  */
  assign n15276_o = yromdo[4];
  /* clock_functions_pack.vhd:101:25  */
  assign n15281_o = c2d10[1];
  /* clock_functions_pack.vhd:101:16  */
  assign n15282_o = n15276_o & n15281_o;
  /* vlm5030_gl.vhd:1691:47  */
  assign n15284_o = xromdo[7];
  /* vlm5030_gl.vhd:1691:37  */
  assign n15285_o = ~n15284_o;
  /* vlm5030_gl.vhd:1691:33  */
  assign n15286_o = tstend2ie | n15285_o;
  /* clock_functions_pack.vhd:147:24  */
  assign n15291_o = nc2d10[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n15292_o = n15286_o | n15291_o;
  /* vlm5030_gl.vhd:1691:18  */
  assign n15293_o = ~n15292_o;
  assign n15295_o = osc[0];
  /* vlm5030_gl.vhd:1697:16  */
  assign n15297_o = {1'b0, mem_block_a};  //  uext
  /* vlm5030_gl.vhd:1697:16  */
  assign n15299_o = $signed(n15297_o) <= $signed(32'b00000000000000000000000000001000);
  /* vlm5030_gl.vhd:1698:18  */
  assign n15300_o = mem_block_a[3:0];  // trunc
  /* vlm5030_gl.vhd:1696:9  */
  assign n15306_o = mem_block_clkmem2 & n15299_o;
  /* vlm5030_gl.vhd:1705:27  */
  assign n15309_o = mem_block_a[3:0];  // trunc
  /* vlm5030_gl.vhd:1705:18  */
  assign n15314_o = ~n20406_data;
  /* vlm5030_gl.vhd:1705:37  */
  assign n15315_o = {1'b0, mem_block_a};  //  uext
  /* vlm5030_gl.vhd:1705:37  */
  assign n15317_o = $signed(n15315_o) <= $signed(32'b00000000000000000000000000001000);
  /* vlm5030_gl.vhd:1705:30  */
  assign n15318_o = n15317_o ? n15314_o : 12'b111111111111;
  assign n15320_o = {n15173_o, n15174_o, n15175_o, n15176_o};
  /* vlm5030_gl.vhd:1715:12  */
  assign arithmetic_block_memxdo = n18906_o; // (signal)
  /* vlm5030_gl.vhd:1716:12  */
  assign arithmetic_block_wl = n15330_o; // (signal)
  /* vlm5030_gl.vhd:1729:12  */
  assign arithmetic_block_row0 = n18910_o; // (signal)
  /* vlm5030_gl.vhd:1729:18  */
  assign arithmetic_block_row1 = n18911_o; // (signal)
  /* vlm5030_gl.vhd:1729:24  */
  assign arithmetic_block_row2 = n18912_o; // (signal)
  /* vlm5030_gl.vhd:1729:30  */
  assign arithmetic_block_row3 = n18913_o; // (signal)
  /* vlm5030_gl.vhd:1729:36  */
  assign arithmetic_block_row4 = n18914_o; // (signal)
  /* vlm5030_gl.vhd:1803:12  */
  assign arithmetic_block_memlatmuxq = n18918_q; // (signal)
  /* vlm5030_gl.vhd:1808:12  */
  assign arithmetic_block_memlatmux = n18919_o; // (signal)
  /* vlm5030_gl.vhd:1816:12  */
  assign arithmetic_block_iereg = n18956_o; // (signal)
  /* vlm5030_gl.vhd:1820:17  */
  assign n15327_o = yromdo[4];
  /* vlm5030_gl.vhd:1820:33  */
  assign n15328_o = yromdo[4];
  /* vlm5030_gl.vhd:1820:23  */
  assign n15329_o = ~n15328_o;
  /* vlm5030_gl.vhd:1820:21  */
  assign n15330_o = {n15327_o, n15329_o};
  /* vlm5030_gl.vhd:1822:40  */
  assign n15332_o = mem1do2ie[11];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15333_o = mem2do2ie[11];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15334_o = {n15332_o, n15333_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15340_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15341_o = n15334_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15342_o = n15340_o & n15341_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15344_o = 1'b0 | n15342_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15346_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15347_o = n15334_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15348_o = n15346_o & n15347_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15349_o = n15344_o | n15348_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15350_o = ~n15349_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15352_o = mem1do2ie[10];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15353_o = mem2do2ie[10];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15354_o = {n15352_o, n15353_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15360_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15361_o = n15354_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15362_o = n15360_o & n15361_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15364_o = 1'b0 | n15362_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15366_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15367_o = n15354_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15368_o = n15366_o & n15367_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15369_o = n15364_o | n15368_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15370_o = ~n15369_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15372_o = mem1do2ie[9];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15373_o = mem2do2ie[9];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15374_o = {n15372_o, n15373_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15380_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15381_o = n15374_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15382_o = n15380_o & n15381_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15384_o = 1'b0 | n15382_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15386_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15387_o = n15374_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15388_o = n15386_o & n15387_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15389_o = n15384_o | n15388_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15390_o = ~n15389_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15392_o = mem1do2ie[8];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15393_o = mem2do2ie[8];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15394_o = {n15392_o, n15393_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15400_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15401_o = n15394_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15402_o = n15400_o & n15401_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15404_o = 1'b0 | n15402_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15406_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15407_o = n15394_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15408_o = n15406_o & n15407_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15409_o = n15404_o | n15408_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15410_o = ~n15409_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15412_o = mem1do2ie[7];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15413_o = mem2do2ie[7];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15414_o = {n15412_o, n15413_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15420_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15421_o = n15414_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15422_o = n15420_o & n15421_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15424_o = 1'b0 | n15422_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15426_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15427_o = n15414_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15428_o = n15426_o & n15427_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15429_o = n15424_o | n15428_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15430_o = ~n15429_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15432_o = mem1do2ie[6];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15433_o = mem2do2ie[6];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15434_o = {n15432_o, n15433_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15440_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15441_o = n15434_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15442_o = n15440_o & n15441_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15444_o = 1'b0 | n15442_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15446_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15447_o = n15434_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15448_o = n15446_o & n15447_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15449_o = n15444_o | n15448_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15450_o = ~n15449_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15452_o = mem1do2ie[5];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15453_o = mem2do2ie[5];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15454_o = {n15452_o, n15453_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15460_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15461_o = n15454_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15462_o = n15460_o & n15461_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15464_o = 1'b0 | n15462_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15466_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15467_o = n15454_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15468_o = n15466_o & n15467_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15469_o = n15464_o | n15468_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15470_o = ~n15469_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15472_o = mem1do2ie[4];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15473_o = mem2do2ie[4];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15474_o = {n15472_o, n15473_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15480_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15481_o = n15474_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15482_o = n15480_o & n15481_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15484_o = 1'b0 | n15482_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15486_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15487_o = n15474_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15488_o = n15486_o & n15487_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15489_o = n15484_o | n15488_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15490_o = ~n15489_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15492_o = mem1do2ie[3];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15493_o = mem2do2ie[3];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15494_o = {n15492_o, n15493_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15500_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15501_o = n15494_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15502_o = n15500_o & n15501_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15504_o = 1'b0 | n15502_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15506_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15507_o = n15494_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15508_o = n15506_o & n15507_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15509_o = n15504_o | n15508_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15510_o = ~n15509_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15512_o = mem1do2ie[2];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15513_o = mem2do2ie[2];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15514_o = {n15512_o, n15513_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15520_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15521_o = n15514_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15522_o = n15520_o & n15521_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15524_o = 1'b0 | n15522_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15526_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15527_o = n15514_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15528_o = n15526_o & n15527_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15529_o = n15524_o | n15528_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15530_o = ~n15529_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15532_o = mem1do2ie[1];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15533_o = mem2do2ie[1];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15534_o = {n15532_o, n15533_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15540_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15541_o = n15534_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15542_o = n15540_o & n15541_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15544_o = 1'b0 | n15542_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15546_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15547_o = n15534_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15548_o = n15546_o & n15547_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15549_o = n15544_o | n15548_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15550_o = ~n15549_o;
  /* vlm5030_gl.vhd:1822:40  */
  assign n15552_o = mem1do2ie[0];
  /* vlm5030_gl.vhd:1822:57  */
  assign n15553_o = mem2do2ie[0];
  /* vlm5030_gl.vhd:1822:46  */
  assign n15554_o = {n15552_o, n15553_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n15560_o = arithmetic_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n15561_o = n15554_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n15562_o = n15560_o & n15561_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15564_o = 1'b0 | n15562_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n15566_o = arithmetic_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n15567_o = n15554_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n15568_o = n15566_o & n15567_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n15569_o = n15564_o | n15568_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n15570_o = ~n15569_o;
  /* vlm5030_gl.vhd:1830:45  */
  assign n15572_o = mem0do[0];
  /* vlm5030_gl.vhd:1752:33  */
  assign n15577_o = ~n15572_o;
  /* vlm5030_gl.vhd:1752:28  */
  assign n15579_o = 1'b1 ^ n15577_o;
  /* vlm5030_gl.vhd:1752:14  */
  assign n15580_o = ~n15579_o;
  /* vlm5030_gl.vhd:1831:30  */
  assign n15581_o = mem0do[0];
  /* vlm5030_gl.vhd:1831:20  */
  assign n15582_o = ~n15581_o;
  /* vlm5030_gl.vhd:1831:45  */
  assign n15583_o = mem0do[1];
  /* vlm5030_gl.vhd:1831:35  */
  assign n15584_o = ~(n15582_o | n15583_o);
  /* vlm5030_gl.vhd:1832:25  */
  assign n15585_o = mem0do[1];
  /* vlm5030_gl.vhd:1833:36  */
  assign n15586_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1838:42  */
  assign n15589_o = arithmetic_block_memxdo[9];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15590_o = ~n15589_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15592_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15593_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15594_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15595_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15596_o = arithmetic_block_row0[3];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15601_o = n15592_o & n15594_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15602_o = n15596_o & n15593_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15603_o = n15601_o | n15602_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15604_o = ~n15603_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15605_o = n15595_o ^ n15604_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15607_o = arithmetic_block_row0[17];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15613_o = n15607_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15615_o = n15613_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15618_o = arithmetic_block_memxdo[8];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15619_o = ~n15618_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15621_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15622_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15623_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15624_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15625_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15630_o = n15621_o & n15623_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15631_o = n15625_o & n15622_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15632_o = n15630_o | n15631_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15633_o = ~n15632_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15634_o = n15624_o ^ n15633_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15636_o = arithmetic_block_row0[18];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15642_o = n15636_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15644_o = n15642_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15647_o = arithmetic_block_memxdo[7];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15648_o = ~n15647_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15650_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15651_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15652_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15653_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15654_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15659_o = n15650_o & n15652_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15660_o = n15654_o & n15651_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15661_o = n15659_o | n15660_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15662_o = ~n15661_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15663_o = n15653_o ^ n15662_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15665_o = arithmetic_block_row0[19];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15671_o = n15665_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15673_o = n15671_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15676_o = arithmetic_block_memxdo[6];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15677_o = ~n15676_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15679_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15680_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15681_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15682_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15683_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15688_o = n15679_o & n15681_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15689_o = n15683_o & n15680_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15690_o = n15688_o | n15689_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15691_o = ~n15690_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15692_o = n15682_o ^ n15691_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15694_o = arithmetic_block_row0[20];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15700_o = n15694_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15702_o = n15700_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15705_o = arithmetic_block_memxdo[5];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15706_o = ~n15705_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15708_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15709_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15710_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15711_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15712_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15717_o = n15708_o & n15710_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15718_o = n15712_o & n15709_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15719_o = n15717_o | n15718_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15720_o = ~n15719_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15721_o = n15711_o ^ n15720_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15723_o = arithmetic_block_row0[21];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15729_o = n15723_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15731_o = n15729_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15734_o = arithmetic_block_memxdo[4];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15735_o = ~n15734_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15737_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15738_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15739_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15740_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15741_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15746_o = n15737_o & n15739_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15747_o = n15741_o & n15738_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15748_o = n15746_o | n15747_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15749_o = ~n15748_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15750_o = n15740_o ^ n15749_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15752_o = arithmetic_block_row0[22];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15758_o = n15752_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15760_o = n15758_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15763_o = arithmetic_block_memxdo[3];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15764_o = ~n15763_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15766_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15767_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15768_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15769_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15770_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15775_o = n15766_o & n15768_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15776_o = n15770_o & n15767_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15777_o = n15775_o | n15776_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15778_o = ~n15777_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15779_o = n15769_o ^ n15778_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15781_o = arithmetic_block_row0[23];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15787_o = n15781_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15789_o = n15787_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15792_o = arithmetic_block_memxdo[2];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15793_o = ~n15792_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15795_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15796_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15797_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15798_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15799_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15804_o = n15795_o & n15797_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15805_o = n15799_o & n15796_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15806_o = n15804_o | n15805_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15807_o = ~n15806_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15808_o = n15798_o ^ n15807_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15810_o = arithmetic_block_row0[24];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15816_o = n15810_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15818_o = n15816_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15821_o = arithmetic_block_memxdo[1];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15822_o = ~n15821_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15824_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15825_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15826_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15827_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15828_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15833_o = n15824_o & n15826_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15834_o = n15828_o & n15825_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15835_o = n15833_o | n15834_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15836_o = ~n15835_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15837_o = n15827_o ^ n15836_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15839_o = arithmetic_block_row0[25];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15845_o = n15839_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15847_o = n15845_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15850_o = arithmetic_block_memxdo[0];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15851_o = ~n15850_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15853_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15854_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15855_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15856_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15857_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15862_o = n15853_o & n15855_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15863_o = n15857_o & n15854_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15864_o = n15862_o | n15863_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15865_o = ~n15864_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15866_o = n15856_o ^ n15865_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15868_o = arithmetic_block_row0[26];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15874_o = n15868_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15876_o = n15874_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15879_o = arithmetic_block_memxdo[11];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15880_o = ~n15879_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15882_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15883_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15884_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15885_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15886_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15891_o = n15882_o & n15884_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15892_o = n15886_o & n15883_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15893_o = n15891_o | n15892_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15894_o = ~n15893_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15895_o = n15885_o ^ n15894_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15897_o = arithmetic_block_row0[27];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15903_o = n15897_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15905_o = n15903_o ^ 1'b0;
  /* vlm5030_gl.vhd:1838:42  */
  assign n15908_o = arithmetic_block_memxdo[10];
  /* vlm5030_gl.vhd:1838:32  */
  assign n15909_o = ~n15908_o;
  /* vlm5030_gl.vhd:1839:61  */
  assign n15911_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1840:48  */
  assign n15912_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1841:48  */
  assign n15913_o = arithmetic_block_row0[1];
  /* vlm5030_gl.vhd:1842:48  */
  assign n15914_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1843:61  */
  assign n15915_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15920_o = n15911_o & n15913_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15921_o = n15915_o & n15912_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15922_o = n15920_o | n15921_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15923_o = ~n15922_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15924_o = n15914_o ^ n15923_o;
  /* vlm5030_gl.vhd:1844:52  */
  assign n15926_o = arithmetic_block_row0[28];
  /* vlm5030_gl.vhd:1783:20  */
  assign n15932_o = n15926_o ^ 1'b0;
  /* vlm5030_gl.vhd:1783:30  */
  assign n15934_o = n15932_o ^ 1'b0;
  /* vlm5030_gl.vhd:1851:34  */
  assign n15936_o = arithmetic_block_row0[0];
  /* vlm5030_gl.vhd:1851:56  */
  assign n15937_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1851:40  */
  assign n15938_o = n15936_o & n15937_o;
  /* vlm5030_gl.vhd:1851:71  */
  assign n15939_o = arithmetic_block_row0[2];
  /* vlm5030_gl.vhd:1851:93  */
  assign n15940_o = arithmetic_block_row0[41];
  /* vlm5030_gl.vhd:1851:81  */
  assign n15941_o = ~n15940_o;
  /* vlm5030_gl.vhd:1851:77  */
  assign n15942_o = n15939_o | n15941_o;
  /* vlm5030_gl.vhd:1851:62  */
  assign n15943_o = n15938_o | n15942_o;
  /* vlm5030_gl.vhd:1851:23  */
  assign n15944_o = ~n15943_o;
  /* vlm5030_gl.vhd:1852:28  */
  assign n15945_o = arithmetic_block_row0[56];
  /* vlm5030_gl.vhd:1857:45  */
  assign n15947_o = mem0do[1];
  /* vlm5030_gl.vhd:1858:45  */
  assign n15948_o = mem0do[2];
  /* vlm5030_gl.vhd:1752:33  */
  assign n15953_o = ~n15948_o;
  /* vlm5030_gl.vhd:1752:28  */
  assign n15954_o = n15947_o ^ n15953_o;
  /* vlm5030_gl.vhd:1752:14  */
  assign n15955_o = ~n15954_o;
  /* vlm5030_gl.vhd:1859:45  */
  assign n15957_o = mem0do[1];
  /* vlm5030_gl.vhd:1860:45  */
  assign n15958_o = mem0do[2];
  /* vlm5030_gl.vhd:1861:45  */
  assign n15959_o = mem0do[3];
  /* vlm5030_gl.vhd:1760:22  */
  assign n15964_o = ~n15957_o;
  /* vlm5030_gl.vhd:1761:22  */
  assign n15965_o = ~n15958_o;
  /* vlm5030_gl.vhd:1761:17  */
  assign n15966_o = n15964_o & n15965_o;
  /* vlm5030_gl.vhd:1762:17  */
  assign n15967_o = n15966_o & n15959_o;
  /* vlm5030_gl.vhd:1765:17  */
  assign n15968_o = n15957_o & n15958_o;
  /* vlm5030_gl.vhd:1766:22  */
  assign n15969_o = ~n15959_o;
  /* vlm5030_gl.vhd:1766:17  */
  assign n15970_o = n15968_o & n15969_o;
  /* vlm5030_gl.vhd:1763:17  */
  assign n15971_o = n15967_o | n15970_o;
  /* vlm5030_gl.vhd:1862:25  */
  assign n15972_o = mem0do[3];
  /* vlm5030_gl.vhd:1866:61  */
  assign n15975_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1867:48  */
  assign n15976_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1868:48  */
  assign n15977_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1869:48  */
  assign n15978_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1870:61  */
  assign n15979_o = arithmetic_block_row0[3];
  /* vlm5030_gl.vhd:1776:41  */
  assign n15984_o = n15975_o & n15977_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n15985_o = n15979_o & n15976_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n15986_o = n15984_o | n15985_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n15987_o = ~n15986_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n15988_o = n15978_o ^ n15987_o;
  /* vlm5030_gl.vhd:1871:41  */
  assign n15989_o = arithmetic_block_row1[17];
  /* vlm5030_gl.vhd:1871:28  */
  assign n15990_o = ~n15989_o;
  /* vlm5030_gl.vhd:1872:32  */
  assign n15993_o = 1'b1 ? 1'b0 : n15994_o;
  /* vlm5030_gl.vhd:1873:38  */
  assign n15994_o = arithmetic_block_row1[17];
  /* vlm5030_gl.vhd:1866:61  */
  assign n15996_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1867:48  */
  assign n15997_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1868:48  */
  assign n15998_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1869:48  */
  assign n15999_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1870:61  */
  assign n16000_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16005_o = n15996_o & n15998_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16006_o = n16000_o & n15997_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16007_o = n16005_o | n16006_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16008_o = ~n16007_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16009_o = n15999_o ^ n16008_o;
  /* vlm5030_gl.vhd:1871:41  */
  assign n16010_o = arithmetic_block_row1[18];
  /* vlm5030_gl.vhd:1871:28  */
  assign n16011_o = ~n16010_o;
  /* vlm5030_gl.vhd:1872:32  */
  assign n16014_o = 1'b0 ? 1'b0 : n16015_o;
  /* vlm5030_gl.vhd:1873:38  */
  assign n16015_o = arithmetic_block_row1[18];
  /* vlm5030_gl.vhd:1876:55  */
  assign n16017_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1877:42  */
  assign n16018_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1878:42  */
  assign n16019_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1879:42  */
  assign n16020_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1880:55  */
  assign n16021_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16026_o = n16017_o & n16019_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16027_o = n16021_o & n16018_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16028_o = n16026_o | n16027_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16029_o = ~n16028_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16030_o = n16020_o ^ n16029_o;
  /* vlm5030_gl.vhd:1881:46  */
  assign n16032_o = arithmetic_block_row1[19];
  /* vlm5030_gl.vhd:1882:45  */
  assign n16033_o = arithmetic_block_row0[30];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16038_o = n16032_o ^ n16033_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16040_o = n16038_o ^ 1'b0;
  /* vlm5030_gl.vhd:1884:36  */
  assign n16041_o = arithmetic_block_row1[19];
  /* vlm5030_gl.vhd:1884:23  */
  assign n16042_o = ~n16041_o;
  /* vlm5030_gl.vhd:1884:54  */
  assign n16043_o = arithmetic_block_row0[30];
  /* vlm5030_gl.vhd:1884:41  */
  assign n16044_o = ~(n16042_o & n16043_o);
  /* vlm5030_gl.vhd:1887:60  */
  assign n16046_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16047_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16048_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16049_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16050_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16055_o = n16046_o & n16048_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16056_o = n16050_o & n16047_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16057_o = n16055_o | n16056_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16058_o = ~n16057_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16059_o = n16049_o ^ n16058_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16061_o = arithmetic_block_row1[20];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16062_o = arithmetic_block_row0[31];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16067_o = n16061_o ^ n16062_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16069_o = n16067_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16071_o = arithmetic_block_row1[20];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16072_o = arithmetic_block_row0[31];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16077_o = n16071_o | n16072_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16079_o = 1'b0 & n16077_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16080_o = n16071_o & n16072_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16081_o = n16079_o | n16080_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16083_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16084_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16085_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16086_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16087_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16092_o = n16083_o & n16085_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16093_o = n16087_o & n16084_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16094_o = n16092_o | n16093_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16095_o = ~n16094_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16096_o = n16086_o ^ n16095_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16098_o = arithmetic_block_row1[21];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16099_o = arithmetic_block_row0[32];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16104_o = n16098_o ^ n16099_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16106_o = n16104_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16108_o = arithmetic_block_row1[21];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16109_o = arithmetic_block_row0[32];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16114_o = n16108_o | n16109_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16116_o = 1'b0 & n16114_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16117_o = n16108_o & n16109_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16118_o = n16116_o | n16117_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16120_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16121_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16122_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16123_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16124_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16129_o = n16120_o & n16122_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16130_o = n16124_o & n16121_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16131_o = n16129_o | n16130_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16132_o = ~n16131_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16133_o = n16123_o ^ n16132_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16135_o = arithmetic_block_row1[22];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16136_o = arithmetic_block_row0[33];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16141_o = n16135_o ^ n16136_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16143_o = n16141_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16145_o = arithmetic_block_row1[22];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16146_o = arithmetic_block_row0[33];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16151_o = n16145_o | n16146_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16153_o = 1'b0 & n16151_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16154_o = n16145_o & n16146_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16155_o = n16153_o | n16154_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16157_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16158_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16159_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16160_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16161_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16166_o = n16157_o & n16159_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16167_o = n16161_o & n16158_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16168_o = n16166_o | n16167_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16169_o = ~n16168_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16170_o = n16160_o ^ n16169_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16172_o = arithmetic_block_row1[23];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16173_o = arithmetic_block_row0[34];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16178_o = n16172_o ^ n16173_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16180_o = n16178_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16182_o = arithmetic_block_row1[23];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16183_o = arithmetic_block_row0[34];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16188_o = n16182_o | n16183_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16190_o = 1'b0 & n16188_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16191_o = n16182_o & n16183_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16192_o = n16190_o | n16191_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16194_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16195_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16196_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16197_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16198_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16203_o = n16194_o & n16196_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16204_o = n16198_o & n16195_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16205_o = n16203_o | n16204_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16206_o = ~n16205_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16207_o = n16197_o ^ n16206_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16209_o = arithmetic_block_row1[24];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16210_o = arithmetic_block_row0[35];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16215_o = n16209_o ^ n16210_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16217_o = n16215_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16219_o = arithmetic_block_row1[24];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16220_o = arithmetic_block_row0[35];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16225_o = n16219_o | n16220_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16227_o = 1'b0 & n16225_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16228_o = n16219_o & n16220_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16229_o = n16227_o | n16228_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16231_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16232_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16233_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16234_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16235_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16240_o = n16231_o & n16233_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16241_o = n16235_o & n16232_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16242_o = n16240_o | n16241_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16243_o = ~n16242_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16244_o = n16234_o ^ n16243_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16246_o = arithmetic_block_row1[25];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16247_o = arithmetic_block_row0[36];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16252_o = n16246_o ^ n16247_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16254_o = n16252_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16256_o = arithmetic_block_row1[25];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16257_o = arithmetic_block_row0[36];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16262_o = n16256_o | n16257_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16264_o = 1'b0 & n16262_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16265_o = n16256_o & n16257_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16266_o = n16264_o | n16265_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16268_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16269_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16270_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16271_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16272_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16277_o = n16268_o & n16270_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16278_o = n16272_o & n16269_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16279_o = n16277_o | n16278_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16280_o = ~n16279_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16281_o = n16271_o ^ n16280_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16283_o = arithmetic_block_row1[26];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16284_o = arithmetic_block_row0[37];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16289_o = n16283_o ^ n16284_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16291_o = n16289_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16293_o = arithmetic_block_row1[26];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16294_o = arithmetic_block_row0[37];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16299_o = n16293_o | n16294_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16301_o = 1'b0 & n16299_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16302_o = n16293_o & n16294_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16303_o = n16301_o | n16302_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16305_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16306_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16307_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16308_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16309_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16314_o = n16305_o & n16307_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16315_o = n16309_o & n16306_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16316_o = n16314_o | n16315_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16317_o = ~n16316_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16318_o = n16308_o ^ n16317_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16320_o = arithmetic_block_row1[27];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16321_o = arithmetic_block_row0[38];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16326_o = n16320_o ^ n16321_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16328_o = n16326_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16330_o = arithmetic_block_row1[27];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16331_o = arithmetic_block_row0[38];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16336_o = n16330_o | n16331_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16338_o = 1'b0 & n16336_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16339_o = n16330_o & n16331_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16340_o = n16338_o | n16339_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16342_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16343_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16344_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16345_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16346_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16351_o = n16342_o & n16344_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16352_o = n16346_o & n16343_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16353_o = n16351_o | n16352_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16354_o = ~n16353_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16355_o = n16345_o ^ n16354_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16357_o = arithmetic_block_row1[28];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16358_o = arithmetic_block_row0[39];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16363_o = n16357_o ^ n16358_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16365_o = n16363_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16367_o = arithmetic_block_row1[28];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16368_o = arithmetic_block_row0[39];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16373_o = n16367_o | n16368_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16375_o = 1'b0 & n16373_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16376_o = n16367_o & n16368_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16377_o = n16375_o | n16376_o;
  /* vlm5030_gl.vhd:1887:60  */
  assign n16379_o = arithmetic_block_row0[16];
  /* vlm5030_gl.vhd:1888:47  */
  assign n16380_o = arithmetic_block_row1[0];
  /* vlm5030_gl.vhd:1889:47  */
  assign n16381_o = arithmetic_block_row1[1];
  /* vlm5030_gl.vhd:1890:47  */
  assign n16382_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1891:60  */
  assign n16383_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16388_o = n16379_o & n16381_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16389_o = n16383_o & n16380_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16390_o = n16388_o | n16389_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16391_o = ~n16390_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16392_o = n16382_o ^ n16391_o;
  /* vlm5030_gl.vhd:1892:52  */
  assign n16394_o = arithmetic_block_row1[29];
  /* vlm5030_gl.vhd:1893:51  */
  assign n16395_o = arithmetic_block_row0[40];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16400_o = n16394_o ^ n16395_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16402_o = n16400_o ^ 1'b0;
  /* vlm5030_gl.vhd:1895:54  */
  assign n16404_o = arithmetic_block_row1[29];
  /* vlm5030_gl.vhd:1896:53  */
  assign n16405_o = arithmetic_block_row0[40];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16410_o = n16404_o | n16405_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16412_o = 1'b0 & n16410_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16413_o = n16404_o & n16405_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16414_o = n16412_o | n16413_o;
  /* vlm5030_gl.vhd:1901:49  */
  assign n16416_o = arithmetic_block_row1[2];
  /* vlm5030_gl.vhd:1901:40  */
  assign n16417_o = ~n16416_o;
  /* vlm5030_gl.vhd:1902:48  */
  assign n16418_o = arithmetic_block_row1[42];
  /* vlm5030_gl.vhd:1903:45  */
  assign n16419_o = arithmetic_block_row0[57];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16424_o = n16417_o | n16418_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16425_o = n16419_o & n16424_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16426_o = n16417_o & n16418_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16427_o = n16425_o | n16426_o;
  /* vlm5030_gl.vhd:1904:50  */
  assign n16429_o = arithmetic_block_row1[55];
  /* vlm5030_gl.vhd:1905:48  */
  assign n16430_o = arithmetic_block_row1[41];
  /* vlm5030_gl.vhd:1906:45  */
  assign n16431_o = arithmetic_block_row1[56];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16436_o = n16429_o | n16430_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16437_o = n16431_o & n16436_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16438_o = n16429_o & n16430_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16439_o = n16437_o | n16438_o;
  /* vlm5030_gl.vhd:1912:45  */
  assign n16441_o = mem0do[3];
  /* vlm5030_gl.vhd:1913:45  */
  assign n16442_o = mem0do[4];
  /* vlm5030_gl.vhd:1752:33  */
  assign n16447_o = ~n16442_o;
  /* vlm5030_gl.vhd:1752:28  */
  assign n16448_o = n16441_o ^ n16447_o;
  /* vlm5030_gl.vhd:1752:14  */
  assign n16449_o = ~n16448_o;
  /* vlm5030_gl.vhd:1914:45  */
  assign n16451_o = mem0do[3];
  /* vlm5030_gl.vhd:1915:45  */
  assign n16452_o = mem0do[4];
  /* vlm5030_gl.vhd:1916:45  */
  assign n16453_o = mem0do[5];
  /* vlm5030_gl.vhd:1760:22  */
  assign n16458_o = ~n16451_o;
  /* vlm5030_gl.vhd:1761:22  */
  assign n16459_o = ~n16452_o;
  /* vlm5030_gl.vhd:1761:17  */
  assign n16460_o = n16458_o & n16459_o;
  /* vlm5030_gl.vhd:1762:17  */
  assign n16461_o = n16460_o & n16453_o;
  /* vlm5030_gl.vhd:1765:17  */
  assign n16462_o = n16451_o & n16452_o;
  /* vlm5030_gl.vhd:1766:22  */
  assign n16463_o = ~n16453_o;
  /* vlm5030_gl.vhd:1766:17  */
  assign n16464_o = n16462_o & n16463_o;
  /* vlm5030_gl.vhd:1763:17  */
  assign n16465_o = n16461_o | n16464_o;
  /* vlm5030_gl.vhd:1917:25  */
  assign n16466_o = mem0do[5];
  /* vlm5030_gl.vhd:1921:61  */
  assign n16469_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1922:48  */
  assign n16470_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1923:48  */
  assign n16471_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1924:48  */
  assign n16472_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1925:61  */
  assign n16473_o = arithmetic_block_row0[3];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16478_o = n16469_o & n16471_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16479_o = n16473_o & n16470_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16480_o = n16478_o | n16479_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16481_o = ~n16480_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16482_o = n16472_o ^ n16481_o;
  /* vlm5030_gl.vhd:1926:41  */
  assign n16483_o = arithmetic_block_row2[17];
  /* vlm5030_gl.vhd:1926:28  */
  assign n16484_o = ~n16483_o;
  /* vlm5030_gl.vhd:1927:32  */
  assign n16487_o = 1'b1 ? 1'b0 : n16488_o;
  /* vlm5030_gl.vhd:1928:38  */
  assign n16488_o = arithmetic_block_row2[17];
  /* vlm5030_gl.vhd:1921:61  */
  assign n16490_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1922:48  */
  assign n16491_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1923:48  */
  assign n16492_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1924:48  */
  assign n16493_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1925:61  */
  assign n16494_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16499_o = n16490_o & n16492_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16500_o = n16494_o & n16491_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16501_o = n16499_o | n16500_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16502_o = ~n16501_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16503_o = n16493_o ^ n16502_o;
  /* vlm5030_gl.vhd:1926:41  */
  assign n16504_o = arithmetic_block_row2[18];
  /* vlm5030_gl.vhd:1926:28  */
  assign n16505_o = ~n16504_o;
  /* vlm5030_gl.vhd:1927:32  */
  assign n16508_o = 1'b0 ? 1'b0 : n16509_o;
  /* vlm5030_gl.vhd:1928:38  */
  assign n16509_o = arithmetic_block_row2[18];
  /* vlm5030_gl.vhd:1932:60  */
  assign n16511_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16512_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16513_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16514_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16515_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16520_o = n16511_o & n16513_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16521_o = n16515_o & n16512_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16522_o = n16520_o | n16521_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16523_o = ~n16522_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16524_o = n16514_o ^ n16523_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16526_o = arithmetic_block_row2[19];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16527_o = arithmetic_block_row1[30];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16528_o = arithmetic_block_row1[44];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16533_o = n16526_o ^ n16527_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16534_o = n16533_o ^ n16528_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16536_o = arithmetic_block_row2[19];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16537_o = arithmetic_block_row1[30];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16538_o = arithmetic_block_row1[44];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16543_o = n16536_o | n16537_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16544_o = n16538_o & n16543_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16545_o = n16536_o & n16537_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16546_o = n16544_o | n16545_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16548_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16549_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16550_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16551_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16552_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16557_o = n16548_o & n16550_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16558_o = n16552_o & n16549_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16559_o = n16557_o | n16558_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16560_o = ~n16559_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16561_o = n16551_o ^ n16560_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16563_o = arithmetic_block_row2[20];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16564_o = arithmetic_block_row1[31];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16565_o = arithmetic_block_row1[45];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16570_o = n16563_o ^ n16564_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16571_o = n16570_o ^ n16565_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16573_o = arithmetic_block_row2[20];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16574_o = arithmetic_block_row1[31];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16575_o = arithmetic_block_row1[45];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16580_o = n16573_o | n16574_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16581_o = n16575_o & n16580_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16582_o = n16573_o & n16574_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16583_o = n16581_o | n16582_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16585_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16586_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16587_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16588_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16589_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16594_o = n16585_o & n16587_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16595_o = n16589_o & n16586_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16596_o = n16594_o | n16595_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16597_o = ~n16596_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16598_o = n16588_o ^ n16597_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16600_o = arithmetic_block_row2[21];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16601_o = arithmetic_block_row1[32];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16602_o = arithmetic_block_row1[46];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16607_o = n16600_o ^ n16601_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16608_o = n16607_o ^ n16602_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16610_o = arithmetic_block_row2[21];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16611_o = arithmetic_block_row1[32];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16612_o = arithmetic_block_row1[46];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16617_o = n16610_o | n16611_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16618_o = n16612_o & n16617_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16619_o = n16610_o & n16611_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16620_o = n16618_o | n16619_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16622_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16623_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16624_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16625_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16626_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16631_o = n16622_o & n16624_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16632_o = n16626_o & n16623_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16633_o = n16631_o | n16632_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16634_o = ~n16633_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16635_o = n16625_o ^ n16634_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16637_o = arithmetic_block_row2[22];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16638_o = arithmetic_block_row1[33];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16639_o = arithmetic_block_row1[47];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16644_o = n16637_o ^ n16638_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16645_o = n16644_o ^ n16639_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16647_o = arithmetic_block_row2[22];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16648_o = arithmetic_block_row1[33];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16649_o = arithmetic_block_row1[47];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16654_o = n16647_o | n16648_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16655_o = n16649_o & n16654_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16656_o = n16647_o & n16648_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16657_o = n16655_o | n16656_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16659_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16660_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16661_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16662_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16663_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16668_o = n16659_o & n16661_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16669_o = n16663_o & n16660_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16670_o = n16668_o | n16669_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16671_o = ~n16670_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16672_o = n16662_o ^ n16671_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16674_o = arithmetic_block_row2[23];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16675_o = arithmetic_block_row1[34];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16676_o = arithmetic_block_row1[48];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16681_o = n16674_o ^ n16675_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16682_o = n16681_o ^ n16676_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16684_o = arithmetic_block_row2[23];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16685_o = arithmetic_block_row1[34];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16686_o = arithmetic_block_row1[48];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16691_o = n16684_o | n16685_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16692_o = n16686_o & n16691_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16693_o = n16684_o & n16685_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16694_o = n16692_o | n16693_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16696_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16697_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16698_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16699_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16700_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16705_o = n16696_o & n16698_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16706_o = n16700_o & n16697_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16707_o = n16705_o | n16706_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16708_o = ~n16707_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16709_o = n16699_o ^ n16708_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16711_o = arithmetic_block_row2[24];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16712_o = arithmetic_block_row1[35];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16713_o = arithmetic_block_row1[49];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16718_o = n16711_o ^ n16712_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16719_o = n16718_o ^ n16713_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16721_o = arithmetic_block_row2[24];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16722_o = arithmetic_block_row1[35];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16723_o = arithmetic_block_row1[49];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16728_o = n16721_o | n16722_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16729_o = n16723_o & n16728_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16730_o = n16721_o & n16722_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16731_o = n16729_o | n16730_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16733_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16734_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16735_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16736_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16737_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16742_o = n16733_o & n16735_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16743_o = n16737_o & n16734_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16744_o = n16742_o | n16743_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16745_o = ~n16744_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16746_o = n16736_o ^ n16745_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16748_o = arithmetic_block_row2[25];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16749_o = arithmetic_block_row1[36];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16750_o = arithmetic_block_row1[50];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16755_o = n16748_o ^ n16749_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16756_o = n16755_o ^ n16750_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16758_o = arithmetic_block_row2[25];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16759_o = arithmetic_block_row1[36];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16760_o = arithmetic_block_row1[50];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16765_o = n16758_o | n16759_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16766_o = n16760_o & n16765_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16767_o = n16758_o & n16759_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16768_o = n16766_o | n16767_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16770_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16771_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16772_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16773_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16774_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16779_o = n16770_o & n16772_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16780_o = n16774_o & n16771_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16781_o = n16779_o | n16780_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16782_o = ~n16781_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16783_o = n16773_o ^ n16782_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16785_o = arithmetic_block_row2[26];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16786_o = arithmetic_block_row1[37];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16787_o = arithmetic_block_row1[51];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16792_o = n16785_o ^ n16786_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16793_o = n16792_o ^ n16787_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16795_o = arithmetic_block_row2[26];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16796_o = arithmetic_block_row1[37];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16797_o = arithmetic_block_row1[51];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16802_o = n16795_o | n16796_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16803_o = n16797_o & n16802_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16804_o = n16795_o & n16796_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16805_o = n16803_o | n16804_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16807_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16808_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16809_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16810_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16811_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16816_o = n16807_o & n16809_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16817_o = n16811_o & n16808_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16818_o = n16816_o | n16817_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16819_o = ~n16818_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16820_o = n16810_o ^ n16819_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16822_o = arithmetic_block_row2[27];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16823_o = arithmetic_block_row1[38];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16824_o = arithmetic_block_row1[52];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16829_o = n16822_o ^ n16823_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16830_o = n16829_o ^ n16824_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16832_o = arithmetic_block_row2[27];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16833_o = arithmetic_block_row1[38];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16834_o = arithmetic_block_row1[52];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16839_o = n16832_o | n16833_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16840_o = n16834_o & n16839_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16841_o = n16832_o & n16833_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16842_o = n16840_o | n16841_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16844_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16845_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16846_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16847_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16848_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16853_o = n16844_o & n16846_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16854_o = n16848_o & n16845_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16855_o = n16853_o | n16854_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16856_o = ~n16855_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16857_o = n16847_o ^ n16856_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16859_o = arithmetic_block_row2[28];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16860_o = arithmetic_block_row1[39];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16861_o = arithmetic_block_row1[53];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16866_o = n16859_o ^ n16860_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16867_o = n16866_o ^ n16861_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16869_o = arithmetic_block_row2[28];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16870_o = arithmetic_block_row1[39];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16871_o = arithmetic_block_row1[53];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16876_o = n16869_o | n16870_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16877_o = n16871_o & n16876_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16878_o = n16869_o & n16870_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16879_o = n16877_o | n16878_o;
  /* vlm5030_gl.vhd:1932:60  */
  assign n16881_o = arithmetic_block_row0[16];
  /* vlm5030_gl.vhd:1933:47  */
  assign n16882_o = arithmetic_block_row2[0];
  /* vlm5030_gl.vhd:1934:47  */
  assign n16883_o = arithmetic_block_row2[1];
  /* vlm5030_gl.vhd:1935:47  */
  assign n16884_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1936:60  */
  assign n16885_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16890_o = n16881_o & n16883_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16891_o = n16885_o & n16882_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16892_o = n16890_o | n16891_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16893_o = ~n16892_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16894_o = n16884_o ^ n16893_o;
  /* vlm5030_gl.vhd:1937:52  */
  assign n16896_o = arithmetic_block_row2[29];
  /* vlm5030_gl.vhd:1938:51  */
  assign n16897_o = arithmetic_block_row1[40];
  /* vlm5030_gl.vhd:1939:53  */
  assign n16898_o = arithmetic_block_row1[54];
  /* vlm5030_gl.vhd:1783:20  */
  assign n16903_o = n16896_o ^ n16897_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n16904_o = n16903_o ^ n16898_o;
  /* vlm5030_gl.vhd:1940:54  */
  assign n16906_o = arithmetic_block_row2[29];
  /* vlm5030_gl.vhd:1941:53  */
  assign n16907_o = arithmetic_block_row1[40];
  /* vlm5030_gl.vhd:1942:55  */
  assign n16908_o = arithmetic_block_row1[54];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16913_o = n16906_o | n16907_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16914_o = n16908_o & n16913_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16915_o = n16906_o & n16907_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16916_o = n16914_o | n16915_o;
  /* vlm5030_gl.vhd:1946:49  */
  assign n16918_o = arithmetic_block_row2[2];
  /* vlm5030_gl.vhd:1946:40  */
  assign n16919_o = ~n16918_o;
  /* vlm5030_gl.vhd:1947:48  */
  assign n16920_o = arithmetic_block_row2[42];
  /* vlm5030_gl.vhd:1948:45  */
  assign n16921_o = arithmetic_block_row1[57];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16926_o = n16919_o | n16920_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16927_o = n16921_o & n16926_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16928_o = n16919_o & n16920_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16929_o = n16927_o | n16928_o;
  /* vlm5030_gl.vhd:1949:50  */
  assign n16931_o = arithmetic_block_row2[55];
  /* vlm5030_gl.vhd:1950:48  */
  assign n16932_o = arithmetic_block_row2[41];
  /* vlm5030_gl.vhd:1951:45  */
  assign n16933_o = arithmetic_block_row2[56];
  /* vlm5030_gl.vhd:1791:34  */
  assign n16938_o = n16931_o | n16932_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n16939_o = n16933_o & n16938_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n16940_o = n16931_o & n16932_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n16941_o = n16939_o | n16940_o;
  /* vlm5030_gl.vhd:1956:45  */
  assign n16943_o = mem0do[5];
  /* vlm5030_gl.vhd:1957:45  */
  assign n16944_o = mem0do[6];
  /* vlm5030_gl.vhd:1752:33  */
  assign n16949_o = ~n16944_o;
  /* vlm5030_gl.vhd:1752:28  */
  assign n16950_o = n16943_o ^ n16949_o;
  /* vlm5030_gl.vhd:1752:14  */
  assign n16951_o = ~n16950_o;
  /* vlm5030_gl.vhd:1958:45  */
  assign n16953_o = mem0do[5];
  /* vlm5030_gl.vhd:1959:45  */
  assign n16954_o = mem0do[6];
  /* vlm5030_gl.vhd:1960:45  */
  assign n16955_o = mem0do[7];
  /* vlm5030_gl.vhd:1760:22  */
  assign n16960_o = ~n16953_o;
  /* vlm5030_gl.vhd:1761:22  */
  assign n16961_o = ~n16954_o;
  /* vlm5030_gl.vhd:1761:17  */
  assign n16962_o = n16960_o & n16961_o;
  /* vlm5030_gl.vhd:1762:17  */
  assign n16963_o = n16962_o & n16955_o;
  /* vlm5030_gl.vhd:1765:17  */
  assign n16964_o = n16953_o & n16954_o;
  /* vlm5030_gl.vhd:1766:22  */
  assign n16965_o = ~n16955_o;
  /* vlm5030_gl.vhd:1766:17  */
  assign n16966_o = n16964_o & n16965_o;
  /* vlm5030_gl.vhd:1763:17  */
  assign n16967_o = n16963_o | n16966_o;
  /* vlm5030_gl.vhd:1961:25  */
  assign n16968_o = mem0do[7];
  /* vlm5030_gl.vhd:1965:61  */
  assign n16971_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1966:48  */
  assign n16972_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1967:48  */
  assign n16973_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1968:48  */
  assign n16974_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1969:61  */
  assign n16975_o = arithmetic_block_row0[3];
  /* vlm5030_gl.vhd:1776:41  */
  assign n16980_o = n16971_o & n16973_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n16981_o = n16975_o & n16972_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n16982_o = n16980_o | n16981_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n16983_o = ~n16982_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n16984_o = n16974_o ^ n16983_o;
  /* vlm5030_gl.vhd:1970:41  */
  assign n16985_o = arithmetic_block_row3[17];
  /* vlm5030_gl.vhd:1970:28  */
  assign n16986_o = ~n16985_o;
  /* vlm5030_gl.vhd:1971:32  */
  assign n16989_o = 1'b1 ? 1'b0 : n16990_o;
  /* vlm5030_gl.vhd:1972:38  */
  assign n16990_o = arithmetic_block_row3[17];
  /* vlm5030_gl.vhd:1965:61  */
  assign n16992_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1966:48  */
  assign n16993_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1967:48  */
  assign n16994_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1968:48  */
  assign n16995_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1969:61  */
  assign n16996_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17001_o = n16992_o & n16994_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17002_o = n16996_o & n16993_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17003_o = n17001_o | n17002_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17004_o = ~n17003_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17005_o = n16995_o ^ n17004_o;
  /* vlm5030_gl.vhd:1970:41  */
  assign n17006_o = arithmetic_block_row3[18];
  /* vlm5030_gl.vhd:1970:28  */
  assign n17007_o = ~n17006_o;
  /* vlm5030_gl.vhd:1971:32  */
  assign n17010_o = 1'b0 ? 1'b0 : n17011_o;
  /* vlm5030_gl.vhd:1972:38  */
  assign n17011_o = arithmetic_block_row3[18];
  /* vlm5030_gl.vhd:1976:60  */
  assign n17013_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17014_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17015_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17016_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17017_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17022_o = n17013_o & n17015_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17023_o = n17017_o & n17014_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17024_o = n17022_o | n17023_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17025_o = ~n17024_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17026_o = n17016_o ^ n17025_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17028_o = arithmetic_block_row3[19];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17029_o = arithmetic_block_row2[30];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17030_o = arithmetic_block_row2[44];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17035_o = n17028_o ^ n17029_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17036_o = n17035_o ^ n17030_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17038_o = arithmetic_block_row3[19];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17039_o = arithmetic_block_row2[30];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17040_o = arithmetic_block_row2[44];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17045_o = n17038_o | n17039_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17046_o = n17040_o & n17045_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17047_o = n17038_o & n17039_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17048_o = n17046_o | n17047_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17050_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17051_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17052_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17053_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17054_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17059_o = n17050_o & n17052_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17060_o = n17054_o & n17051_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17061_o = n17059_o | n17060_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17062_o = ~n17061_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17063_o = n17053_o ^ n17062_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17065_o = arithmetic_block_row3[20];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17066_o = arithmetic_block_row2[31];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17067_o = arithmetic_block_row2[45];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17072_o = n17065_o ^ n17066_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17073_o = n17072_o ^ n17067_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17075_o = arithmetic_block_row3[20];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17076_o = arithmetic_block_row2[31];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17077_o = arithmetic_block_row2[45];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17082_o = n17075_o | n17076_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17083_o = n17077_o & n17082_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17084_o = n17075_o & n17076_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17085_o = n17083_o | n17084_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17087_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17088_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17089_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17090_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17091_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17096_o = n17087_o & n17089_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17097_o = n17091_o & n17088_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17098_o = n17096_o | n17097_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17099_o = ~n17098_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17100_o = n17090_o ^ n17099_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17102_o = arithmetic_block_row3[21];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17103_o = arithmetic_block_row2[32];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17104_o = arithmetic_block_row2[46];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17109_o = n17102_o ^ n17103_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17110_o = n17109_o ^ n17104_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17112_o = arithmetic_block_row3[21];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17113_o = arithmetic_block_row2[32];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17114_o = arithmetic_block_row2[46];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17119_o = n17112_o | n17113_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17120_o = n17114_o & n17119_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17121_o = n17112_o & n17113_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17122_o = n17120_o | n17121_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17124_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17125_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17126_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17127_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17128_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17133_o = n17124_o & n17126_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17134_o = n17128_o & n17125_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17135_o = n17133_o | n17134_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17136_o = ~n17135_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17137_o = n17127_o ^ n17136_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17139_o = arithmetic_block_row3[22];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17140_o = arithmetic_block_row2[33];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17141_o = arithmetic_block_row2[47];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17146_o = n17139_o ^ n17140_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17147_o = n17146_o ^ n17141_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17149_o = arithmetic_block_row3[22];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17150_o = arithmetic_block_row2[33];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17151_o = arithmetic_block_row2[47];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17156_o = n17149_o | n17150_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17157_o = n17151_o & n17156_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17158_o = n17149_o & n17150_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17159_o = n17157_o | n17158_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17161_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17162_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17163_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17164_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17165_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17170_o = n17161_o & n17163_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17171_o = n17165_o & n17162_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17172_o = n17170_o | n17171_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17173_o = ~n17172_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17174_o = n17164_o ^ n17173_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17176_o = arithmetic_block_row3[23];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17177_o = arithmetic_block_row2[34];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17178_o = arithmetic_block_row2[48];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17183_o = n17176_o ^ n17177_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17184_o = n17183_o ^ n17178_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17186_o = arithmetic_block_row3[23];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17187_o = arithmetic_block_row2[34];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17188_o = arithmetic_block_row2[48];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17193_o = n17186_o | n17187_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17194_o = n17188_o & n17193_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17195_o = n17186_o & n17187_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17196_o = n17194_o | n17195_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17198_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17199_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17200_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17201_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17202_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17207_o = n17198_o & n17200_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17208_o = n17202_o & n17199_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17209_o = n17207_o | n17208_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17210_o = ~n17209_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17211_o = n17201_o ^ n17210_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17213_o = arithmetic_block_row3[24];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17214_o = arithmetic_block_row2[35];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17215_o = arithmetic_block_row2[49];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17220_o = n17213_o ^ n17214_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17221_o = n17220_o ^ n17215_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17223_o = arithmetic_block_row3[24];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17224_o = arithmetic_block_row2[35];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17225_o = arithmetic_block_row2[49];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17230_o = n17223_o | n17224_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17231_o = n17225_o & n17230_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17232_o = n17223_o & n17224_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17233_o = n17231_o | n17232_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17235_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17236_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17237_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17238_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17239_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17244_o = n17235_o & n17237_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17245_o = n17239_o & n17236_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17246_o = n17244_o | n17245_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17247_o = ~n17246_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17248_o = n17238_o ^ n17247_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17250_o = arithmetic_block_row3[25];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17251_o = arithmetic_block_row2[36];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17252_o = arithmetic_block_row2[50];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17257_o = n17250_o ^ n17251_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17258_o = n17257_o ^ n17252_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17260_o = arithmetic_block_row3[25];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17261_o = arithmetic_block_row2[36];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17262_o = arithmetic_block_row2[50];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17267_o = n17260_o | n17261_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17268_o = n17262_o & n17267_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17269_o = n17260_o & n17261_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17270_o = n17268_o | n17269_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17272_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17273_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17274_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17275_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17276_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17281_o = n17272_o & n17274_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17282_o = n17276_o & n17273_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17283_o = n17281_o | n17282_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17284_o = ~n17283_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17285_o = n17275_o ^ n17284_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17287_o = arithmetic_block_row3[26];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17288_o = arithmetic_block_row2[37];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17289_o = arithmetic_block_row2[51];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17294_o = n17287_o ^ n17288_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17295_o = n17294_o ^ n17289_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17297_o = arithmetic_block_row3[26];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17298_o = arithmetic_block_row2[37];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17299_o = arithmetic_block_row2[51];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17304_o = n17297_o | n17298_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17305_o = n17299_o & n17304_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17306_o = n17297_o & n17298_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17307_o = n17305_o | n17306_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17309_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17310_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17311_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17312_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17313_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17318_o = n17309_o & n17311_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17319_o = n17313_o & n17310_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17320_o = n17318_o | n17319_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17321_o = ~n17320_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17322_o = n17312_o ^ n17321_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17324_o = arithmetic_block_row3[27];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17325_o = arithmetic_block_row2[38];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17326_o = arithmetic_block_row2[52];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17331_o = n17324_o ^ n17325_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17332_o = n17331_o ^ n17326_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17334_o = arithmetic_block_row3[27];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17335_o = arithmetic_block_row2[38];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17336_o = arithmetic_block_row2[52];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17341_o = n17334_o | n17335_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17342_o = n17336_o & n17341_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17343_o = n17334_o & n17335_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17344_o = n17342_o | n17343_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17346_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17347_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17348_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17349_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17350_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17355_o = n17346_o & n17348_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17356_o = n17350_o & n17347_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17357_o = n17355_o | n17356_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17358_o = ~n17357_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17359_o = n17349_o ^ n17358_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17361_o = arithmetic_block_row3[28];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17362_o = arithmetic_block_row2[39];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17363_o = arithmetic_block_row2[53];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17368_o = n17361_o ^ n17362_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17369_o = n17368_o ^ n17363_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17371_o = arithmetic_block_row3[28];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17372_o = arithmetic_block_row2[39];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17373_o = arithmetic_block_row2[53];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17378_o = n17371_o | n17372_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17379_o = n17373_o & n17378_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17380_o = n17371_o & n17372_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17381_o = n17379_o | n17380_o;
  /* vlm5030_gl.vhd:1976:60  */
  assign n17383_o = arithmetic_block_row0[16];
  /* vlm5030_gl.vhd:1977:47  */
  assign n17384_o = arithmetic_block_row3[0];
  /* vlm5030_gl.vhd:1978:47  */
  assign n17385_o = arithmetic_block_row3[1];
  /* vlm5030_gl.vhd:1979:47  */
  assign n17386_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1980:60  */
  assign n17387_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17392_o = n17383_o & n17385_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17393_o = n17387_o & n17384_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17394_o = n17392_o | n17393_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17395_o = ~n17394_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17396_o = n17386_o ^ n17395_o;
  /* vlm5030_gl.vhd:1981:52  */
  assign n17398_o = arithmetic_block_row3[29];
  /* vlm5030_gl.vhd:1982:51  */
  assign n17399_o = arithmetic_block_row2[40];
  /* vlm5030_gl.vhd:1983:53  */
  assign n17400_o = arithmetic_block_row2[54];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17405_o = n17398_o ^ n17399_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17406_o = n17405_o ^ n17400_o;
  /* vlm5030_gl.vhd:1984:54  */
  assign n17408_o = arithmetic_block_row3[29];
  /* vlm5030_gl.vhd:1985:53  */
  assign n17409_o = arithmetic_block_row2[40];
  /* vlm5030_gl.vhd:1986:55  */
  assign n17410_o = arithmetic_block_row2[54];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17415_o = n17408_o | n17409_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17416_o = n17410_o & n17415_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17417_o = n17408_o & n17409_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17418_o = n17416_o | n17417_o;
  /* vlm5030_gl.vhd:1990:49  */
  assign n17420_o = arithmetic_block_row3[2];
  /* vlm5030_gl.vhd:1990:40  */
  assign n17421_o = ~n17420_o;
  /* vlm5030_gl.vhd:1991:48  */
  assign n17422_o = arithmetic_block_row3[42];
  /* vlm5030_gl.vhd:1992:45  */
  assign n17423_o = arithmetic_block_row2[57];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17428_o = n17421_o | n17422_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17429_o = n17423_o & n17428_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17430_o = n17421_o & n17422_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17431_o = n17429_o | n17430_o;
  /* vlm5030_gl.vhd:1993:50  */
  assign n17433_o = arithmetic_block_row3[55];
  /* vlm5030_gl.vhd:1994:48  */
  assign n17434_o = arithmetic_block_row3[41];
  /* vlm5030_gl.vhd:1995:45  */
  assign n17435_o = arithmetic_block_row3[56];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17440_o = n17433_o | n17434_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17441_o = n17435_o & n17440_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17442_o = n17433_o & n17434_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17443_o = n17441_o | n17442_o;
  /* vlm5030_gl.vhd:2000:45  */
  assign n17445_o = mem0do[7];
  /* vlm5030_gl.vhd:2001:45  */
  assign n17446_o = mem0do[8];
  /* vlm5030_gl.vhd:1752:33  */
  assign n17451_o = ~n17446_o;
  /* vlm5030_gl.vhd:1752:28  */
  assign n17452_o = n17445_o ^ n17451_o;
  /* vlm5030_gl.vhd:1752:14  */
  assign n17453_o = ~n17452_o;
  /* vlm5030_gl.vhd:2002:45  */
  assign n17455_o = mem0do[7];
  /* vlm5030_gl.vhd:2003:45  */
  assign n17456_o = mem0do[8];
  /* vlm5030_gl.vhd:2004:45  */
  assign n17457_o = mem0do[9];
  /* vlm5030_gl.vhd:1760:22  */
  assign n17462_o = ~n17455_o;
  /* vlm5030_gl.vhd:1761:22  */
  assign n17463_o = ~n17456_o;
  /* vlm5030_gl.vhd:1761:17  */
  assign n17464_o = n17462_o & n17463_o;
  /* vlm5030_gl.vhd:1762:17  */
  assign n17465_o = n17464_o & n17457_o;
  /* vlm5030_gl.vhd:1765:17  */
  assign n17466_o = n17455_o & n17456_o;
  /* vlm5030_gl.vhd:1766:22  */
  assign n17467_o = ~n17457_o;
  /* vlm5030_gl.vhd:1766:17  */
  assign n17468_o = n17466_o & n17467_o;
  /* vlm5030_gl.vhd:1763:17  */
  assign n17469_o = n17465_o | n17468_o;
  /* vlm5030_gl.vhd:2005:25  */
  assign n17470_o = mem0do[9];
  /* vlm5030_gl.vhd:2009:61  */
  assign n17473_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:2010:48  */
  assign n17474_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2011:48  */
  assign n17475_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2012:48  */
  assign n17476_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2013:61  */
  assign n17477_o = arithmetic_block_row0[3];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17482_o = n17473_o & n17475_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17483_o = n17477_o & n17474_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17484_o = n17482_o | n17483_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17485_o = ~n17484_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17486_o = n17476_o ^ n17485_o;
  /* vlm5030_gl.vhd:2014:41  */
  assign n17487_o = arithmetic_block_row4[17];
  /* vlm5030_gl.vhd:2014:28  */
  assign n17488_o = ~n17487_o;
  /* vlm5030_gl.vhd:2015:32  */
  assign n17491_o = 1'b1 ? 1'b0 : n17492_o;
  /* vlm5030_gl.vhd:2016:38  */
  assign n17492_o = arithmetic_block_row4[17];
  /* vlm5030_gl.vhd:2009:61  */
  assign n17494_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:2010:48  */
  assign n17495_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2011:48  */
  assign n17496_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2012:48  */
  assign n17497_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2013:61  */
  assign n17498_o = arithmetic_block_row0[4];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17503_o = n17494_o & n17496_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17504_o = n17498_o & n17495_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17505_o = n17503_o | n17504_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17506_o = ~n17505_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17507_o = n17497_o ^ n17506_o;
  /* vlm5030_gl.vhd:2014:41  */
  assign n17508_o = arithmetic_block_row4[18];
  /* vlm5030_gl.vhd:2014:28  */
  assign n17509_o = ~n17508_o;
  /* vlm5030_gl.vhd:2015:32  */
  assign n17512_o = 1'b0 ? 1'b0 : n17513_o;
  /* vlm5030_gl.vhd:2016:38  */
  assign n17513_o = arithmetic_block_row4[18];
  /* vlm5030_gl.vhd:2020:60  */
  assign n17515_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17516_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17517_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17518_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17519_o = arithmetic_block_row0[5];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17524_o = n17515_o & n17517_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17525_o = n17519_o & n17516_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17526_o = n17524_o | n17525_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17527_o = ~n17526_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17528_o = n17518_o ^ n17527_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17530_o = arithmetic_block_row4[19];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17531_o = arithmetic_block_row3[30];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17532_o = arithmetic_block_row3[44];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17537_o = n17530_o ^ n17531_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17538_o = n17537_o ^ n17532_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17540_o = arithmetic_block_row4[19];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17541_o = arithmetic_block_row3[30];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17542_o = arithmetic_block_row3[44];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17547_o = n17540_o | n17541_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17548_o = n17542_o & n17547_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17549_o = n17540_o & n17541_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17550_o = n17548_o | n17549_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17552_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17553_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17554_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17555_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17556_o = arithmetic_block_row0[6];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17561_o = n17552_o & n17554_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17562_o = n17556_o & n17553_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17563_o = n17561_o | n17562_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17564_o = ~n17563_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17565_o = n17555_o ^ n17564_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17567_o = arithmetic_block_row4[20];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17568_o = arithmetic_block_row3[31];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17569_o = arithmetic_block_row3[45];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17574_o = n17567_o ^ n17568_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17575_o = n17574_o ^ n17569_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17577_o = arithmetic_block_row4[20];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17578_o = arithmetic_block_row3[31];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17579_o = arithmetic_block_row3[45];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17584_o = n17577_o | n17578_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17585_o = n17579_o & n17584_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17586_o = n17577_o & n17578_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17587_o = n17585_o | n17586_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17589_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17590_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17591_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17592_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17593_o = arithmetic_block_row0[7];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17598_o = n17589_o & n17591_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17599_o = n17593_o & n17590_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17600_o = n17598_o | n17599_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17601_o = ~n17600_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17602_o = n17592_o ^ n17601_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17604_o = arithmetic_block_row4[21];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17605_o = arithmetic_block_row3[32];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17606_o = arithmetic_block_row3[46];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17611_o = n17604_o ^ n17605_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17612_o = n17611_o ^ n17606_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17614_o = arithmetic_block_row4[21];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17615_o = arithmetic_block_row3[32];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17616_o = arithmetic_block_row3[46];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17621_o = n17614_o | n17615_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17622_o = n17616_o & n17621_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17623_o = n17614_o & n17615_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17624_o = n17622_o | n17623_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17626_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17627_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17628_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17629_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17630_o = arithmetic_block_row0[8];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17635_o = n17626_o & n17628_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17636_o = n17630_o & n17627_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17637_o = n17635_o | n17636_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17638_o = ~n17637_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17639_o = n17629_o ^ n17638_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17641_o = arithmetic_block_row4[22];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17642_o = arithmetic_block_row3[33];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17643_o = arithmetic_block_row3[47];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17648_o = n17641_o ^ n17642_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17649_o = n17648_o ^ n17643_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17651_o = arithmetic_block_row4[22];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17652_o = arithmetic_block_row3[33];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17653_o = arithmetic_block_row3[47];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17658_o = n17651_o | n17652_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17659_o = n17653_o & n17658_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17660_o = n17651_o & n17652_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17661_o = n17659_o | n17660_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17663_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17664_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17665_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17666_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17667_o = arithmetic_block_row0[9];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17672_o = n17663_o & n17665_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17673_o = n17667_o & n17664_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17674_o = n17672_o | n17673_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17675_o = ~n17674_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17676_o = n17666_o ^ n17675_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17678_o = arithmetic_block_row4[23];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17679_o = arithmetic_block_row3[34];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17680_o = arithmetic_block_row3[48];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17685_o = n17678_o ^ n17679_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17686_o = n17685_o ^ n17680_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17688_o = arithmetic_block_row4[23];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17689_o = arithmetic_block_row3[34];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17690_o = arithmetic_block_row3[48];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17695_o = n17688_o | n17689_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17696_o = n17690_o & n17695_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17697_o = n17688_o & n17689_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17698_o = n17696_o | n17697_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17700_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17701_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17702_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17703_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17704_o = arithmetic_block_row0[10];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17709_o = n17700_o & n17702_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17710_o = n17704_o & n17701_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17711_o = n17709_o | n17710_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17712_o = ~n17711_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17713_o = n17703_o ^ n17712_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17715_o = arithmetic_block_row4[24];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17716_o = arithmetic_block_row3[35];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17717_o = arithmetic_block_row3[49];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17722_o = n17715_o ^ n17716_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17723_o = n17722_o ^ n17717_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17725_o = arithmetic_block_row4[24];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17726_o = arithmetic_block_row3[35];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17727_o = arithmetic_block_row3[49];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17732_o = n17725_o | n17726_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17733_o = n17727_o & n17732_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17734_o = n17725_o & n17726_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17735_o = n17733_o | n17734_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17737_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17738_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17739_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17740_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17741_o = arithmetic_block_row0[11];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17746_o = n17737_o & n17739_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17747_o = n17741_o & n17738_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17748_o = n17746_o | n17747_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17749_o = ~n17748_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17750_o = n17740_o ^ n17749_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17752_o = arithmetic_block_row4[25];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17753_o = arithmetic_block_row3[36];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17754_o = arithmetic_block_row3[50];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17759_o = n17752_o ^ n17753_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17760_o = n17759_o ^ n17754_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17762_o = arithmetic_block_row4[25];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17763_o = arithmetic_block_row3[36];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17764_o = arithmetic_block_row3[50];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17769_o = n17762_o | n17763_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17770_o = n17764_o & n17769_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17771_o = n17762_o & n17763_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17772_o = n17770_o | n17771_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17774_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17775_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17776_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17777_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17778_o = arithmetic_block_row0[12];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17783_o = n17774_o & n17776_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17784_o = n17778_o & n17775_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17785_o = n17783_o | n17784_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17786_o = ~n17785_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17787_o = n17777_o ^ n17786_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17789_o = arithmetic_block_row4[26];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17790_o = arithmetic_block_row3[37];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17791_o = arithmetic_block_row3[51];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17796_o = n17789_o ^ n17790_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17797_o = n17796_o ^ n17791_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17799_o = arithmetic_block_row4[26];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17800_o = arithmetic_block_row3[37];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17801_o = arithmetic_block_row3[51];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17806_o = n17799_o | n17800_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17807_o = n17801_o & n17806_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17808_o = n17799_o & n17800_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17809_o = n17807_o | n17808_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17811_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17812_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17813_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17814_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17815_o = arithmetic_block_row0[13];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17820_o = n17811_o & n17813_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17821_o = n17815_o & n17812_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17822_o = n17820_o | n17821_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17823_o = ~n17822_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17824_o = n17814_o ^ n17823_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17826_o = arithmetic_block_row4[27];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17827_o = arithmetic_block_row3[38];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17828_o = arithmetic_block_row3[52];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17833_o = n17826_o ^ n17827_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17834_o = n17833_o ^ n17828_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17836_o = arithmetic_block_row4[27];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17837_o = arithmetic_block_row3[38];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17838_o = arithmetic_block_row3[52];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17843_o = n17836_o | n17837_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17844_o = n17838_o & n17843_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17845_o = n17836_o & n17837_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17846_o = n17844_o | n17845_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17848_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17849_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17850_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17851_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17852_o = arithmetic_block_row0[14];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17857_o = n17848_o & n17850_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17858_o = n17852_o & n17849_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17859_o = n17857_o | n17858_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17860_o = ~n17859_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17861_o = n17851_o ^ n17860_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17863_o = arithmetic_block_row4[28];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17864_o = arithmetic_block_row3[39];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17865_o = arithmetic_block_row3[53];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17870_o = n17863_o ^ n17864_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17871_o = n17870_o ^ n17865_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17873_o = arithmetic_block_row4[28];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17874_o = arithmetic_block_row3[39];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17875_o = arithmetic_block_row3[53];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17880_o = n17873_o | n17874_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17881_o = n17875_o & n17880_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17882_o = n17873_o & n17874_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17883_o = n17881_o | n17882_o;
  /* vlm5030_gl.vhd:2020:60  */
  assign n17885_o = arithmetic_block_row0[16];
  /* vlm5030_gl.vhd:2021:47  */
  assign n17886_o = arithmetic_block_row4[0];
  /* vlm5030_gl.vhd:2022:47  */
  assign n17887_o = arithmetic_block_row4[1];
  /* vlm5030_gl.vhd:2023:47  */
  assign n17888_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2024:60  */
  assign n17889_o = arithmetic_block_row0[15];
  /* vlm5030_gl.vhd:1776:41  */
  assign n17894_o = n17885_o & n17887_o;
  /* vlm5030_gl.vhd:1776:68  */
  assign n17895_o = n17889_o & n17886_o;
  /* vlm5030_gl.vhd:1776:52  */
  assign n17896_o = n17894_o | n17895_o;
  /* vlm5030_gl.vhd:1776:24  */
  assign n17897_o = ~n17896_o;
  /* vlm5030_gl.vhd:1776:20  */
  assign n17898_o = n17888_o ^ n17897_o;
  /* vlm5030_gl.vhd:2025:52  */
  assign n17900_o = arithmetic_block_row4[29];
  /* vlm5030_gl.vhd:2026:51  */
  assign n17901_o = arithmetic_block_row3[40];
  /* vlm5030_gl.vhd:2027:53  */
  assign n17902_o = arithmetic_block_row3[54];
  /* vlm5030_gl.vhd:1783:20  */
  assign n17907_o = n17900_o ^ n17901_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n17908_o = n17907_o ^ n17902_o;
  /* vlm5030_gl.vhd:2028:54  */
  assign n17910_o = arithmetic_block_row4[29];
  /* vlm5030_gl.vhd:2029:53  */
  assign n17911_o = arithmetic_block_row3[40];
  /* vlm5030_gl.vhd:2030:55  */
  assign n17912_o = arithmetic_block_row3[54];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17917_o = n17910_o | n17911_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17918_o = n17912_o & n17917_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17919_o = n17910_o & n17911_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17920_o = n17918_o | n17919_o;
  /* vlm5030_gl.vhd:2034:49  */
  assign n17922_o = arithmetic_block_row4[2];
  /* vlm5030_gl.vhd:2034:40  */
  assign n17923_o = ~n17922_o;
  /* vlm5030_gl.vhd:2035:48  */
  assign n17924_o = arithmetic_block_row4[42];
  /* vlm5030_gl.vhd:2036:45  */
  assign n17925_o = arithmetic_block_row3[57];
  /* vlm5030_gl.vhd:1791:34  */
  assign n17930_o = n17923_o | n17924_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n17931_o = n17925_o & n17930_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n17932_o = n17923_o & n17924_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n17933_o = n17931_o | n17932_o;
  /* vlm5030_gl.vhd:2037:28  */
  assign n17934_o = arithmetic_block_row4[56];
  assign n17941_o = c2d7fin[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n17943_o = c2d7fin[2];
  /* vlm5030_gl.vhd:2046:23  */
  assign n17945_o = ~ieregdrv;
  /* vlm5030_gl.vhd:2051:45  */
  assign n17948_o = arithmetic_block_row4[44];
  /* clock_functions_pack.vhd:175:17  */
  assign n17954_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n17955_o = ~n17954_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n17956_o = n17955_o ? n17948_o : n17960_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n17957_o = arithmetic_block_memlatmuxq[0];
  /* vlm5030_gl.vhd:2052:66  */
  assign n17958_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n17959_o = ~n17958_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n17960_o = n17959_o ? n17957_o : n17962_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n17961_o = arithmetic_block_memlatmuxq[0];
  /* vlm5030_gl.vhd:2053:31  */
  assign n17962_o = ~n17961_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n17963_o = arithmetic_block_row4[30];
  /* vlm5030_gl.vhd:2051:45  */
  assign n17964_o = arithmetic_block_row4[45];
  /* clock_functions_pack.vhd:175:17  */
  assign n17970_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n17971_o = ~n17970_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n17972_o = n17971_o ? n17964_o : n17976_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n17973_o = arithmetic_block_memlatmuxq[1];
  /* vlm5030_gl.vhd:2052:66  */
  assign n17974_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n17975_o = ~n17974_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n17976_o = n17975_o ? n17973_o : n17978_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n17977_o = arithmetic_block_memlatmuxq[1];
  /* vlm5030_gl.vhd:2053:31  */
  assign n17978_o = ~n17977_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n17979_o = arithmetic_block_row4[31];
  /* vlm5030_gl.vhd:2051:45  */
  assign n17980_o = arithmetic_block_row4[46];
  /* clock_functions_pack.vhd:175:17  */
  assign n17986_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n17987_o = ~n17986_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n17988_o = n17987_o ? n17980_o : n17992_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n17989_o = arithmetic_block_memlatmuxq[2];
  /* vlm5030_gl.vhd:2052:66  */
  assign n17990_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n17991_o = ~n17990_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n17992_o = n17991_o ? n17989_o : n17994_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n17993_o = arithmetic_block_memlatmuxq[2];
  /* vlm5030_gl.vhd:2053:31  */
  assign n17994_o = ~n17993_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n17995_o = arithmetic_block_row4[32];
  /* vlm5030_gl.vhd:2051:45  */
  assign n17996_o = arithmetic_block_row4[47];
  /* clock_functions_pack.vhd:175:17  */
  assign n18002_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18003_o = ~n18002_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18004_o = n18003_o ? n17996_o : n18008_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18005_o = arithmetic_block_memlatmuxq[3];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18006_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18007_o = ~n18006_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18008_o = n18007_o ? n18005_o : n18010_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18009_o = arithmetic_block_memlatmuxq[3];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18010_o = ~n18009_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18011_o = arithmetic_block_row4[33];
  /* vlm5030_gl.vhd:2051:45  */
  assign n18012_o = arithmetic_block_row4[48];
  /* clock_functions_pack.vhd:175:17  */
  assign n18018_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18019_o = ~n18018_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18020_o = n18019_o ? n18012_o : n18024_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18021_o = arithmetic_block_memlatmuxq[4];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18022_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18023_o = ~n18022_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18024_o = n18023_o ? n18021_o : n18026_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18025_o = arithmetic_block_memlatmuxq[4];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18026_o = ~n18025_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18027_o = arithmetic_block_row4[34];
  /* vlm5030_gl.vhd:2051:45  */
  assign n18028_o = arithmetic_block_row4[49];
  /* clock_functions_pack.vhd:175:17  */
  assign n18034_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18035_o = ~n18034_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18036_o = n18035_o ? n18028_o : n18040_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18037_o = arithmetic_block_memlatmuxq[5];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18038_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18039_o = ~n18038_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18040_o = n18039_o ? n18037_o : n18042_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18041_o = arithmetic_block_memlatmuxq[5];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18042_o = ~n18041_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18043_o = arithmetic_block_row4[35];
  /* vlm5030_gl.vhd:2051:45  */
  assign n18044_o = arithmetic_block_row4[50];
  /* clock_functions_pack.vhd:175:17  */
  assign n18050_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18051_o = ~n18050_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18052_o = n18051_o ? n18044_o : n18056_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18053_o = arithmetic_block_memlatmuxq[6];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18054_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18055_o = ~n18054_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18056_o = n18055_o ? n18053_o : n18058_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18057_o = arithmetic_block_memlatmuxq[6];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18058_o = ~n18057_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18059_o = arithmetic_block_row4[36];
  /* vlm5030_gl.vhd:2051:45  */
  assign n18060_o = arithmetic_block_row4[51];
  /* clock_functions_pack.vhd:175:17  */
  assign n18066_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18067_o = ~n18066_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18068_o = n18067_o ? n18060_o : n18072_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18069_o = arithmetic_block_memlatmuxq[7];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18070_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18071_o = ~n18070_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18072_o = n18071_o ? n18069_o : n18074_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18073_o = arithmetic_block_memlatmuxq[7];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18074_o = ~n18073_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18075_o = arithmetic_block_row4[37];
  /* vlm5030_gl.vhd:2051:45  */
  assign n18076_o = arithmetic_block_row4[52];
  /* clock_functions_pack.vhd:175:17  */
  assign n18082_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18083_o = ~n18082_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18084_o = n18083_o ? n18076_o : n18088_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18085_o = arithmetic_block_memlatmuxq[8];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18086_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18087_o = ~n18086_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18088_o = n18087_o ? n18085_o : n18090_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18089_o = arithmetic_block_memlatmuxq[8];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18090_o = ~n18089_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18091_o = arithmetic_block_row4[38];
  /* vlm5030_gl.vhd:2051:45  */
  assign n18092_o = arithmetic_block_row4[53];
  /* clock_functions_pack.vhd:175:17  */
  assign n18098_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18099_o = ~n18098_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18100_o = n18099_o ? n18092_o : n18104_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18101_o = arithmetic_block_memlatmuxq[9];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18102_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18103_o = ~n18102_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18104_o = n18103_o ? n18101_o : n18106_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18105_o = arithmetic_block_memlatmuxq[9];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18106_o = ~n18105_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18107_o = arithmetic_block_row4[39];
  /* vlm5030_gl.vhd:2051:45  */
  assign n18108_o = arithmetic_block_row4[54];
  /* clock_functions_pack.vhd:175:17  */
  assign n18114_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18115_o = ~n18114_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18116_o = n18115_o ? n18108_o : n18120_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18117_o = arithmetic_block_memlatmuxq[10];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18118_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18119_o = ~n18118_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18120_o = n18119_o ? n18117_o : n18122_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18121_o = arithmetic_block_memlatmuxq[10];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18122_o = ~n18121_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18123_o = arithmetic_block_row4[40];
  /* vlm5030_gl.vhd:2051:45  */
  assign n18124_o = arithmetic_block_row4[55];
  /* clock_functions_pack.vhd:175:17  */
  assign n18130_o = c2d7fin[1];
  /* clock_functions_pack.vhd:175:21  */
  assign n18131_o = ~n18130_o;
  /* vlm5030_gl.vhd:2051:55  */
  assign n18132_o = n18131_o ? n18124_o : n18136_o;
  /* vlm5030_gl.vhd:2052:45  */
  assign n18133_o = arithmetic_block_memlatmuxq[11];
  /* vlm5030_gl.vhd:2052:66  */
  assign n18134_o = yromdo[4];
  /* vlm5030_gl.vhd:2052:70  */
  assign n18135_o = ~n18134_o;
  /* vlm5030_gl.vhd:2051:74  */
  assign n18136_o = n18135_o ? n18133_o : n18138_o;
  /* vlm5030_gl.vhd:2053:45  */
  assign n18137_o = arithmetic_block_memlatmuxq[11];
  /* vlm5030_gl.vhd:2053:31  */
  assign n18138_o = ~n18137_o;
  /* vlm5030_gl.vhd:2054:41  */
  assign n18139_o = arithmetic_block_row4[41];
  /* vlm5030_gl.vhd:2063:46  */
  assign n18140_o = yromdo[4];
  /* vlm5030_gl.vhd:2063:36  */
  assign n18141_o = ~n18140_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18147_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2063:50  */
  assign n18148_o = n18147_o ? n18141_o : n18149_o;
  /* vlm5030_gl.vhd:2064:41  */
  assign n18149_o = arithmetic_block_row4[57];
  assign n18156_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18158_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18162_o = nie[9];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18166_o = arithmetic_block_iereg[0];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18167_o = ~n18166_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18173_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18174_o = n18173_o ? n18167_o : n18175_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18175_o = arithmetic_block_memlatmux[12];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18177_o = arithmetic_block_memlatmux[0];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18178_o = arithmetic_block_iereg[12];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18179_o = arithmetic_block_iereg[25];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18184_o = n18177_o | n18178_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18185_o = n18179_o & n18184_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18186_o = n18177_o & n18178_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18187_o = n18185_o | n18186_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18189_o = arithmetic_block_memlatmux[0];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18190_o = arithmetic_block_iereg[12];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18191_o = arithmetic_block_iereg[25];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18196_o = n18189_o ^ n18190_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18197_o = n18196_o ^ n18191_o;
  assign n18204_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18206_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18210_o = nie[8];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18214_o = arithmetic_block_iereg[1];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18215_o = ~n18214_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18221_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18222_o = n18221_o ? n18215_o : n18223_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18223_o = arithmetic_block_memlatmux[13];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18225_o = arithmetic_block_memlatmux[1];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18226_o = arithmetic_block_iereg[13];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18227_o = arithmetic_block_iereg[26];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18232_o = n18225_o | n18226_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18233_o = n18227_o & n18232_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18234_o = n18225_o & n18226_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18235_o = n18233_o | n18234_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18237_o = arithmetic_block_memlatmux[1];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18238_o = arithmetic_block_iereg[13];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18239_o = arithmetic_block_iereg[26];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18244_o = n18237_o ^ n18238_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18245_o = n18244_o ^ n18239_o;
  assign n18252_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18254_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18258_o = nie[7];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18262_o = arithmetic_block_iereg[2];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18263_o = ~n18262_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18269_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18270_o = n18269_o ? n18263_o : n18271_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18271_o = arithmetic_block_memlatmux[14];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18273_o = arithmetic_block_memlatmux[2];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18274_o = arithmetic_block_iereg[14];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18275_o = arithmetic_block_iereg[27];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18280_o = n18273_o | n18274_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18281_o = n18275_o & n18280_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18282_o = n18273_o & n18274_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18283_o = n18281_o | n18282_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18285_o = arithmetic_block_memlatmux[2];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18286_o = arithmetic_block_iereg[14];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18287_o = arithmetic_block_iereg[27];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18292_o = n18285_o ^ n18286_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18293_o = n18292_o ^ n18287_o;
  assign n18300_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18302_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18306_o = nie[6];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18310_o = arithmetic_block_iereg[3];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18311_o = ~n18310_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18317_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18318_o = n18317_o ? n18311_o : n18319_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18319_o = arithmetic_block_memlatmux[15];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18321_o = arithmetic_block_memlatmux[3];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18322_o = arithmetic_block_iereg[15];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18323_o = arithmetic_block_iereg[28];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18328_o = n18321_o | n18322_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18329_o = n18323_o & n18328_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18330_o = n18321_o & n18322_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18331_o = n18329_o | n18330_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18333_o = arithmetic_block_memlatmux[3];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18334_o = arithmetic_block_iereg[15];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18335_o = arithmetic_block_iereg[28];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18340_o = n18333_o ^ n18334_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18341_o = n18340_o ^ n18335_o;
  assign n18348_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18350_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18354_o = nie[5];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18358_o = arithmetic_block_iereg[4];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18359_o = ~n18358_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18365_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18366_o = n18365_o ? n18359_o : n18367_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18367_o = arithmetic_block_memlatmux[16];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18369_o = arithmetic_block_memlatmux[4];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18370_o = arithmetic_block_iereg[16];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18371_o = arithmetic_block_iereg[29];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18376_o = n18369_o | n18370_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18377_o = n18371_o & n18376_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18378_o = n18369_o & n18370_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18379_o = n18377_o | n18378_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18381_o = arithmetic_block_memlatmux[4];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18382_o = arithmetic_block_iereg[16];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18383_o = arithmetic_block_iereg[29];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18388_o = n18381_o ^ n18382_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18389_o = n18388_o ^ n18383_o;
  assign n18396_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18398_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18402_o = nie[4];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18406_o = arithmetic_block_iereg[5];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18407_o = ~n18406_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18413_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18414_o = n18413_o ? n18407_o : n18415_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18415_o = arithmetic_block_memlatmux[17];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18417_o = arithmetic_block_memlatmux[5];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18418_o = arithmetic_block_iereg[17];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18419_o = arithmetic_block_iereg[30];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18424_o = n18417_o | n18418_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18425_o = n18419_o & n18424_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18426_o = n18417_o & n18418_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18427_o = n18425_o | n18426_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18429_o = arithmetic_block_memlatmux[5];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18430_o = arithmetic_block_iereg[17];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18431_o = arithmetic_block_iereg[30];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18436_o = n18429_o ^ n18430_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18437_o = n18436_o ^ n18431_o;
  assign n18444_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18446_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18450_o = nie[3];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18454_o = arithmetic_block_iereg[6];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18455_o = ~n18454_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18461_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18462_o = n18461_o ? n18455_o : n18463_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18463_o = arithmetic_block_memlatmux[18];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18465_o = arithmetic_block_memlatmux[6];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18466_o = arithmetic_block_iereg[18];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18467_o = arithmetic_block_iereg[31];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18472_o = n18465_o | n18466_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18473_o = n18467_o & n18472_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18474_o = n18465_o & n18466_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18475_o = n18473_o | n18474_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18477_o = arithmetic_block_memlatmux[6];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18478_o = arithmetic_block_iereg[18];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18479_o = arithmetic_block_iereg[31];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18484_o = n18477_o ^ n18478_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18485_o = n18484_o ^ n18479_o;
  assign n18492_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18494_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18498_o = nie[2];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18502_o = arithmetic_block_iereg[7];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18503_o = ~n18502_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18509_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18510_o = n18509_o ? n18503_o : n18511_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18511_o = arithmetic_block_memlatmux[19];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18513_o = arithmetic_block_memlatmux[7];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18514_o = arithmetic_block_iereg[19];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18515_o = arithmetic_block_iereg[32];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18520_o = n18513_o | n18514_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18521_o = n18515_o & n18520_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18522_o = n18513_o & n18514_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18523_o = n18521_o | n18522_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18525_o = arithmetic_block_memlatmux[7];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18526_o = arithmetic_block_iereg[19];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18527_o = arithmetic_block_iereg[32];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18532_o = n18525_o ^ n18526_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18533_o = n18532_o ^ n18527_o;
  assign n18540_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18542_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18546_o = nie[1];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18550_o = arithmetic_block_iereg[8];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18551_o = ~n18550_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18557_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18558_o = n18557_o ? n18551_o : n18559_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18559_o = arithmetic_block_memlatmux[20];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18561_o = arithmetic_block_memlatmux[8];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18562_o = arithmetic_block_iereg[20];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18563_o = arithmetic_block_iereg[33];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18568_o = n18561_o | n18562_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18569_o = n18563_o & n18568_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18570_o = n18561_o & n18562_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18571_o = n18569_o | n18570_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18573_o = arithmetic_block_memlatmux[8];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18574_o = arithmetic_block_iereg[20];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18575_o = arithmetic_block_iereg[33];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18580_o = n18573_o ^ n18574_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18581_o = n18580_o ^ n18575_o;
  assign n18588_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18590_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18594_o = nie[0];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18598_o = arithmetic_block_iereg[9];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18599_o = ~n18598_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18605_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18606_o = n18605_o ? n18599_o : n18607_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18607_o = arithmetic_block_memlatmux[21];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18609_o = arithmetic_block_memlatmux[9];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18610_o = arithmetic_block_iereg[21];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18611_o = arithmetic_block_iereg[34];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18616_o = n18609_o | n18610_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18617_o = n18611_o & n18616_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18618_o = n18609_o & n18610_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18619_o = n18617_o | n18618_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18621_o = arithmetic_block_memlatmux[9];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18622_o = arithmetic_block_iereg[21];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18623_o = arithmetic_block_iereg[34];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18628_o = n18621_o ^ n18622_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18629_o = n18628_o ^ n18623_o;
  assign n18636_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18638_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18642_o = nie[11];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18646_o = arithmetic_block_iereg[10];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18647_o = ~n18646_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18653_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18654_o = n18653_o ? n18647_o : n18655_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18655_o = arithmetic_block_memlatmux[22];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18657_o = arithmetic_block_memlatmux[10];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18658_o = arithmetic_block_iereg[22];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18659_o = arithmetic_block_iereg[35];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18664_o = n18657_o | n18658_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18665_o = n18659_o & n18664_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18666_o = n18657_o & n18658_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18667_o = n18665_o | n18666_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18669_o = arithmetic_block_memlatmux[10];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18670_o = arithmetic_block_iereg[22];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18671_o = arithmetic_block_iereg[35];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18676_o = n18669_o ^ n18670_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18677_o = n18676_o ^ n18671_o;
  assign n18684_o = ieregload[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18686_o = ieregload[3];
  /* vlm5030_gl.vhd:2071:32  */
  assign n18690_o = nie[10];
  /* vlm5030_gl.vhd:2075:40  */
  assign n18694_o = arithmetic_block_iereg[11];
  /* vlm5030_gl.vhd:2075:29  */
  assign n18695_o = ~n18694_o;
  /* clock_functions_pack.vhd:175:17  */
  assign n18701_o = c2d7fin[1];
  /* vlm5030_gl.vhd:2075:48  */
  assign n18702_o = n18701_o ? n18695_o : n18703_o;
  /* vlm5030_gl.vhd:2076:44  */
  assign n18703_o = arithmetic_block_memlatmux[23];
  /* vlm5030_gl.vhd:2077:59  */
  assign n18705_o = arithmetic_block_memlatmux[11];
  /* vlm5030_gl.vhd:2078:57  */
  assign n18706_o = arithmetic_block_iereg[23];
  /* vlm5030_gl.vhd:2079:56  */
  assign n18707_o = arithmetic_block_iereg[36];
  /* vlm5030_gl.vhd:1791:34  */
  assign n18712_o = n18705_o | n18706_o;
  /* vlm5030_gl.vhd:1791:23  */
  assign n18713_o = n18707_o & n18712_o;
  /* vlm5030_gl.vhd:1793:23  */
  assign n18714_o = n18705_o & n18706_o;
  /* vlm5030_gl.vhd:1792:17  */
  assign n18715_o = n18713_o | n18714_o;
  /* vlm5030_gl.vhd:2080:57  */
  assign n18717_o = arithmetic_block_memlatmux[11];
  /* vlm5030_gl.vhd:2081:55  */
  assign n18718_o = arithmetic_block_iereg[23];
  /* vlm5030_gl.vhd:2082:54  */
  assign n18719_o = arithmetic_block_iereg[36];
  /* vlm5030_gl.vhd:1783:20  */
  assign n18724_o = n18717_o ^ n18718_o;
  /* vlm5030_gl.vhd:1783:30  */
  assign n18725_o = n18724_o ^ n18719_o;
  /* vlm5030_gl.vhd:2085:23  */
  assign n18726_o = arithmetic_block_iereg[48:37];
  /* vlm5030_gl.vhd:2085:58  */
  assign n18728_o = arithmetic_block_iereg[24];
  /* vlm5030_gl.vhd:2085:44  */
  assign n18729_o = ~n18728_o;
  /* vlm5030_gl.vhd:2085:82  */
  assign n18730_o = arithmetic_block_iereg[25];
  /* vlm5030_gl.vhd:2085:68  */
  assign n18731_o = ~n18730_o;
  /* vlm5030_gl.vhd:2085:63  */
  assign n18732_o = n18729_o ^ n18731_o;
  /* clock_functions_pack.vhd:124:26  */
  assign n18737_o = c2d7fin[1];
  /* clock_functions_pack.vhd:124:16  */
  assign n18738_o = ~(n18732_o & n18737_o);
  /* vlm5030_gl.vhd:2085:33  */
  assign n18739_o = n18738_o ? n18726_o : n18753_o;
  /* vlm5030_gl.vhd:2086:58  */
  assign n18742_o = arithmetic_block_iereg[25];
  /* vlm5030_gl.vhd:2086:82  */
  assign n18743_o = arithmetic_block_iereg[24];
  /* vlm5030_gl.vhd:2086:68  */
  assign n18744_o = ~n18743_o;
  /* vlm5030_gl.vhd:2086:64  */
  assign n18745_o = n18742_o | n18744_o;
  /* clock_functions_pack.vhd:147:24  */
  assign n18750_o = nc2d7fin[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n18751_o = n18745_o | n18750_o;
  /* vlm5030_gl.vhd:2086:38  */
  assign n18752_o = ~n18751_o;
  /* vlm5030_gl.vhd:2085:110  */
  assign n18753_o = n18752_o ? 12'b111111111111 : n18767_o;
  /* vlm5030_gl.vhd:2087:58  */
  assign n18756_o = arithmetic_block_iereg[25];
  /* vlm5030_gl.vhd:2087:44  */
  assign n18757_o = ~n18756_o;
  /* vlm5030_gl.vhd:2087:82  */
  assign n18758_o = arithmetic_block_iereg[24];
  /* vlm5030_gl.vhd:2087:64  */
  assign n18759_o = n18757_o | n18758_o;
  /* clock_functions_pack.vhd:147:24  */
  assign n18764_o = nc2d7fin[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n18765_o = n18759_o | n18764_o;
  /* vlm5030_gl.vhd:2087:38  */
  assign n18766_o = ~n18765_o;
  /* vlm5030_gl.vhd:2086:110  */
  assign n18767_o = n18766_o ? 12'b000000000000 : 12'bX;
  /* vlm5030_gl.vhd:2090:37  */
  assign n18771_o = ieregdrv[9];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18774_o = ieregdrv[8];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18777_o = ieregdrv[7];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18780_o = ieregdrv[6];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18783_o = ieregdrv[5];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18786_o = ieregdrv[4];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18789_o = ieregdrv[3];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18792_o = ieregdrv[2];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18795_o = ieregdrv[1];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18798_o = ieregdrv[0];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18801_o = ieregdrv[11];
  /* vlm5030_gl.vhd:2090:37  */
  assign n18804_o = ieregdrv[10];
  /* vlm5030_gl.vhd:2093:37  */
  assign n18807_o = yromdo[4];
  /* clock_functions_pack.vhd:93:26  */
  assign n18812_o = c2d10[0];
  /* clock_functions_pack.vhd:94:26  */
  assign n18813_o = c2d10[1];
  /* clock_functions_pack.vhd:94:30  */
  assign n18814_o = n18813_o & n18807_o;
  /* clock_functions_pack.vhd:95:26  */
  assign n18815_o = c2d10[2];
  /* clock_functions_pack.vhd:95:31  */
  assign n18816_o = n18815_o & n18807_o;
  /* clock_functions_pack.vhd:96:26  */
  assign n18817_o = c2d10[3];
  /* clock_functions_pack.vhd:96:31  */
  assign n18818_o = n18817_o & n18807_o;
  assign n18819_o = {n18818_o, n18816_o, n18814_o, n18812_o};
  /* vlm5030_gl.vhd:2093:78  */
  assign n18821_o = yromdo[4];
  /* vlm5030_gl.vhd:2093:67  */
  assign n18822_o = ~(xromdo7q & n18821_o);
  /* clock_functions_pack.vhd:93:26  */
  assign n18827_o = c2d6[0];
  /* clock_functions_pack.vhd:94:26  */
  assign n18828_o = c2d6[1];
  /* clock_functions_pack.vhd:94:30  */
  assign n18829_o = n18828_o & n18822_o;
  /* clock_functions_pack.vhd:95:26  */
  assign n18830_o = c2d6[2];
  /* clock_functions_pack.vhd:95:31  */
  assign n18831_o = n18830_o & n18822_o;
  /* clock_functions_pack.vhd:96:26  */
  assign n18832_o = c2d6[3];
  /* clock_functions_pack.vhd:96:31  */
  assign n18833_o = n18832_o & n18822_o;
  assign n18834_o = {n18833_o, n18831_o, n18829_o, n18827_o};
  /* clock_functions_pack.vhd:129:26  */
  assign n18839_o = n18819_o[0];
  /* clock_functions_pack.vhd:130:26  */
  assign n18840_o = n18819_o[1];
  /* clock_functions_pack.vhd:130:38  */
  assign n18841_o = n18834_o[1];
  /* clock_functions_pack.vhd:130:30  */
  assign n18842_o = n18840_o | n18841_o;
  /* clock_functions_pack.vhd:131:27  */
  assign n18843_o = n18819_o[2];
  /* clock_functions_pack.vhd:131:45  */
  assign n18844_o = n18834_o[1];
  /* clock_functions_pack.vhd:131:36  */
  assign n18845_o = ~n18844_o;
  /* clock_functions_pack.vhd:131:32  */
  assign n18846_o = n18843_o & n18845_o;
  /* clock_functions_pack.vhd:132:27  */
  assign n18847_o = n18834_o[2];
  /* clock_functions_pack.vhd:132:45  */
  assign n18848_o = n18819_o[1];
  /* clock_functions_pack.vhd:132:36  */
  assign n18849_o = ~n18848_o;
  /* clock_functions_pack.vhd:132:32  */
  assign n18850_o = n18847_o & n18849_o;
  /* clock_functions_pack.vhd:131:50  */
  assign n18851_o = n18846_o | n18850_o;
  /* clock_functions_pack.vhd:133:27  */
  assign n18852_o = n18819_o[3];
  /* clock_functions_pack.vhd:133:45  */
  assign n18853_o = n18834_o[1];
  /* clock_functions_pack.vhd:133:36  */
  assign n18854_o = ~n18853_o;
  /* clock_functions_pack.vhd:133:32  */
  assign n18855_o = n18852_o & n18854_o;
  /* clock_functions_pack.vhd:133:62  */
  assign n18856_o = n18834_o[2];
  /* clock_functions_pack.vhd:133:53  */
  assign n18857_o = ~n18856_o;
  /* clock_functions_pack.vhd:133:49  */
  assign n18858_o = n18855_o & n18857_o;
  /* clock_functions_pack.vhd:134:27  */
  assign n18859_o = n18834_o[3];
  /* clock_functions_pack.vhd:134:45  */
  assign n18860_o = n18819_o[1];
  /* clock_functions_pack.vhd:134:36  */
  assign n18861_o = ~n18860_o;
  /* clock_functions_pack.vhd:134:32  */
  assign n18862_o = n18859_o & n18861_o;
  /* clock_functions_pack.vhd:134:62  */
  assign n18863_o = n18819_o[2];
  /* clock_functions_pack.vhd:134:53  */
  assign n18864_o = ~n18863_o;
  /* clock_functions_pack.vhd:134:49  */
  assign n18865_o = n18862_o & n18864_o;
  /* clock_functions_pack.vhd:133:68  */
  assign n18866_o = n18858_o | n18865_o;
  assign n18867_o = {n18866_o, n18851_o, n18842_o, n18839_o};
  /* vlm5030_gl.vhd:2094:45  */
  assign n18869_o = xromdo[7];
  /* vlm5030_gl.vhd:2094:36  */
  assign n18870_o = tstend2ie | n18869_o;
  /* clock_functions_pack.vhd:147:24  */
  assign n18875_o = nc2d10[1];
  /* clock_functions_pack.vhd:147:16  */
  assign n18876_o = n18870_o | n18875_o;
  /* vlm5030_gl.vhd:2094:21  */
  assign n18877_o = ~n18876_o;
  /* vlm5030_gl.vhd:2100:33  */
  assign n18879_o = xromdo[9];
  /* clock_functions_pack.vhd:93:26  */
  assign n18884_o = c2d10[0];
  /* clock_functions_pack.vhd:94:26  */
  assign n18885_o = c2d10[1];
  /* clock_functions_pack.vhd:94:30  */
  assign n18886_o = n18885_o & n18879_o;
  /* clock_functions_pack.vhd:95:26  */
  assign n18887_o = c2d10[2];
  /* clock_functions_pack.vhd:95:31  */
  assign n18888_o = n18887_o & n18879_o;
  /* clock_functions_pack.vhd:96:26  */
  assign n18889_o = c2d10[3];
  /* clock_functions_pack.vhd:96:31  */
  assign n18890_o = n18889_o & n18879_o;
  assign n18891_o = {n18890_o, n18888_o, n18886_o, n18884_o};
  /* vlm5030_gl.vhd:2101:22  */
  assign n18892_o = ~(i_tst1 | xromdo7q);
  assign n18899_o = c2d10xr9[0];
  /* clock_functions_pack.vhd:70:42  */
  assign n18901_o = c2d10xr9[3];
  /* vlm5030_gl.vhd:2106:22  */
  assign n18903_o = ~nie;
  assign n18906_o = {n15350_o, n15370_o, n15390_o, n15410_o, n15430_o, n15450_o, n15470_o, n15490_o, n15510_o, n15530_o, n15550_o, n15570_o};
  assign n18910_o = {n15945_o, n15944_o, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n15934_o, n15905_o, n15876_o, n15847_o, n15818_o, n15789_o, n15760_o, n15731_o, n15702_o, n15673_o, n15644_o, n15615_o, 1'b0, n15924_o, n15895_o, n15866_o, n15837_o, n15808_o, n15779_o, n15750_o, n15721_o, n15692_o, n15663_o, n15634_o, n15605_o, 1'b0, n15909_o, n15880_o, n15851_o, n15822_o, n15793_o, n15764_o, n15735_o, n15706_o, n15677_o, n15648_o, n15619_o, n15590_o, n15586_o, n15585_o, n15584_o, n15580_o};
  assign n18911_o = {n16439_o, n16427_o, n16414_o, n16377_o, n16340_o, n16303_o, n16266_o, n16229_o, n16192_o, n16155_o, n16118_o, n16081_o, n16044_o, n16014_o, n15993_o, n16402_o, n16365_o, n16328_o, n16291_o, n16254_o, n16217_o, n16180_o, n16143_o, n16106_o, n16069_o, n16040_o, n16011_o, n15990_o, n16392_o, n16355_o, n16318_o, n16281_o, n16244_o, n16207_o, n16170_o, n16133_o, n16096_o, n16059_o, n16030_o, n16009_o, n15988_o, 14'b00000000000000, n15972_o, n15971_o, n15955_o};
  assign n18912_o = {n16941_o, n16929_o, n16916_o, n16879_o, n16842_o, n16805_o, n16768_o, n16731_o, n16694_o, n16657_o, n16620_o, n16583_o, n16546_o, n16508_o, n16487_o, n16904_o, n16867_o, n16830_o, n16793_o, n16756_o, n16719_o, n16682_o, n16645_o, n16608_o, n16571_o, n16534_o, n16505_o, n16484_o, n16894_o, n16857_o, n16820_o, n16783_o, n16746_o, n16709_o, n16672_o, n16635_o, n16598_o, n16561_o, n16524_o, n16503_o, n16482_o, 14'b00000000000000, n16466_o, n16465_o, n16449_o};
  assign n18913_o = {n17443_o, n17431_o, n17418_o, n17381_o, n17344_o, n17307_o, n17270_o, n17233_o, n17196_o, n17159_o, n17122_o, n17085_o, n17048_o, n17010_o, n16989_o, n17406_o, n17369_o, n17332_o, n17295_o, n17258_o, n17221_o, n17184_o, n17147_o, n17110_o, n17073_o, n17036_o, n17007_o, n16986_o, n17396_o, n17359_o, n17322_o, n17285_o, n17248_o, n17211_o, n17174_o, n17137_o, n17100_o, n17063_o, n17026_o, n17005_o, n16984_o, 14'b00000000000000, n16968_o, n16967_o, n16951_o};
  assign n18914_o = {n17934_o, n17933_o, n17920_o, n17883_o, n17846_o, n17809_o, n17772_o, n17735_o, n17698_o, n17661_o, n17624_o, n17587_o, n17550_o, n17512_o, n17491_o, n17908_o, n17871_o, n17834_o, n17797_o, n17760_o, n17723_o, n17686_o, n17649_o, n17612_o, n17575_o, n17538_o, n17509_o, n17488_o, n17898_o, n17861_o, n17824_o, n17787_o, n17750_o, n17713_o, n17676_o, n17639_o, n17602_o, n17565_o, n17528_o, n17507_o, n17486_o, 14'b00000000000000, n17470_o, n17469_o, n17453_o};
  /* vlm5030_gl.vhd:2045:7  */
  assign n18917_o = n17943_o ? n17945_o : arithmetic_block_memlatmuxq;
  /* vlm5030_gl.vhd:2045:7  */
  always @(posedge n17941_o)
    n18918_q <= n18917_o;
  /* vlm5030_gl.vhd:2045:7  */
  assign n18919_o = {n18139_o, n18123_o, n18107_o, n18091_o, n18075_o, n18059_o, n18043_o, n18027_o, n18011_o, n17995_o, n17979_o, n17963_o, n18132_o, n18116_o, n18100_o, n18084_o, n18068_o, n18052_o, n18036_o, n18020_o, n18004_o, n17988_o, n17972_o, n17956_o};
  assign n18920_o = arithmetic_block_iereg[11];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18921_o = n18686_o ? n18690_o : n18920_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18684_o)
    n18922_q <= n18921_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18923_o = arithmetic_block_iereg[10];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18924_o = n18638_o ? n18642_o : n18923_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18636_o)
    n18925_q <= n18924_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18926_o = arithmetic_block_iereg[9];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18927_o = n18590_o ? n18594_o : n18926_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18588_o)
    n18928_q <= n18927_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18929_o = arithmetic_block_iereg[8];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18930_o = n18542_o ? n18546_o : n18929_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18540_o)
    n18931_q <= n18930_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18932_o = arithmetic_block_iereg[7];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18933_o = n18494_o ? n18498_o : n18932_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18492_o)
    n18934_q <= n18933_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18935_o = arithmetic_block_iereg[6];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18936_o = n18446_o ? n18450_o : n18935_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18444_o)
    n18937_q <= n18936_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18938_o = arithmetic_block_iereg[5];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18939_o = n18398_o ? n18402_o : n18938_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18396_o)
    n18940_q <= n18939_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18941_o = arithmetic_block_iereg[4];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18942_o = n18350_o ? n18354_o : n18941_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18348_o)
    n18943_q <= n18942_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18944_o = arithmetic_block_iereg[3];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18945_o = n18302_o ? n18306_o : n18944_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18300_o)
    n18946_q <= n18945_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18947_o = arithmetic_block_iereg[2];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18948_o = n18254_o ? n18258_o : n18947_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18252_o)
    n18949_q <= n18948_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18950_o = arithmetic_block_iereg[1];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18951_o = n18206_o ? n18210_o : n18950_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18204_o)
    n18952_q <= n18951_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18953_o = arithmetic_block_iereg[0];
  /* vlm5030_gl.vhd:2070:9  */
  assign n18954_o = n18158_o ? n18162_o : n18953_o;
  /* vlm5030_gl.vhd:2070:9  */
  always @(posedge n18156_o)
    n18955_q <= n18954_o;
  /* vlm5030_gl.vhd:2070:9  */
  assign n18956_o = {n18725_o, n18677_o, n18629_o, n18581_o, n18533_o, n18485_o, n18437_o, n18389_o, n18341_o, n18293_o, n18245_o, n18197_o, n18148_o, n18715_o, n18667_o, n18619_o, n18571_o, n18523_o, n18475_o, n18427_o, n18379_o, n18331_o, n18283_o, n18235_o, n18187_o, n18702_o, n18654_o, n18606_o, n18558_o, n18510_o, n18462_o, n18414_o, n18366_o, n18318_o, n18270_o, n18222_o, n18174_o, n18922_q, n18925_q, n18928_q, n18931_q, n18934_q, n18937_q, n18940_q, n18943_q, n18946_q, n18949_q, n18952_q, n18955_q};
  /* vlm5030_gl.vhd:2117:12  */
  assign nie_block_wl = n18961_o; // (signal)
  /* vlm5030_gl.vhd:2120:38  */
  assign n18957_o = {enidlinv2ie, enidl2ie};
  /* vlm5030_gl.vhd:2120:49  */
  assign n18958_o = {n18957_o, enmem12ie};
  /* vlm5030_gl.vhd:2120:65  */
  assign n18959_o = {n18958_o, enmem22ie};
  /* vlm5030_gl.vhd:2120:81  */
  assign n18960_o = {n18959_o, enieregfa2ie};
  /* vlm5030_gl.vhd:2120:99  */
  assign n18961_o = {n18960_o, tstend2ie};
  /* vlm5030_gl.vhd:2122:60  */
  assign n18963_o = mem1do2ie[0];
  /* vlm5030_gl.vhd:2122:49  */
  assign n18965_o = {2'b01, n18963_o};
  /* vlm5030_gl.vhd:2122:76  */
  assign n18966_o = mem2do2ie[0];
  /* vlm5030_gl.vhd:2122:65  */
  assign n18967_o = {n18965_o, n18966_o};
  /* vlm5030_gl.vhd:2122:94  */
  assign n18968_o = ieregdrv4ie[0];
  /* vlm5030_gl.vhd:2122:81  */
  assign n18969_o = {n18967_o, n18968_o};
  /* vlm5030_gl.vhd:2122:105  */
  assign n18970_o = i_d[0];
  /* vlm5030_gl.vhd:2122:99  */
  assign n18971_o = {n18969_o, n18970_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n18977_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n18978_o = n18971_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n18979_o = n18977_o & n18978_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n18981_o = 1'b0 | n18979_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n18983_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n18984_o = n18971_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n18985_o = n18983_o & n18984_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n18986_o = n18981_o | n18985_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n18987_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n18988_o = n18971_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n18989_o = n18987_o & n18988_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n18990_o = n18986_o | n18989_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n18991_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n18992_o = n18971_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n18993_o = n18991_o & n18992_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n18994_o = n18990_o | n18993_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n18995_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n18996_o = n18971_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n18997_o = n18995_o & n18996_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n18998_o = n18994_o | n18997_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n18999_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19000_o = n18971_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19001_o = n18999_o & n19000_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19002_o = n18998_o | n19001_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19003_o = ~n19002_o;
  /* vlm5030_gl.vhd:2123:34  */
  assign n19005_o = idlat[0];
  /* vlm5030_gl.vhd:2123:25  */
  assign n19006_o = ~n19005_o;
  /* vlm5030_gl.vhd:2123:45  */
  assign n19007_o = idlat[0];
  /* vlm5030_gl.vhd:2123:38  */
  assign n19008_o = {n19006_o, n19007_o};
  /* vlm5030_gl.vhd:2123:60  */
  assign n19009_o = mem1do2ie[1];
  /* vlm5030_gl.vhd:2123:49  */
  assign n19010_o = {n19008_o, n19009_o};
  /* vlm5030_gl.vhd:2123:76  */
  assign n19011_o = mem2do2ie[1];
  /* vlm5030_gl.vhd:2123:65  */
  assign n19012_o = {n19010_o, n19011_o};
  /* vlm5030_gl.vhd:2123:94  */
  assign n19013_o = ieregdrv4ie[1];
  /* vlm5030_gl.vhd:2123:81  */
  assign n19014_o = {n19012_o, n19013_o};
  /* vlm5030_gl.vhd:2123:105  */
  assign n19015_o = i_d[1];
  /* vlm5030_gl.vhd:2123:99  */
  assign n19016_o = {n19014_o, n19015_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19022_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19023_o = n19016_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19024_o = n19022_o & n19023_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19026_o = 1'b0 | n19024_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19028_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19029_o = n19016_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19030_o = n19028_o & n19029_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19031_o = n19026_o | n19030_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19032_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19033_o = n19016_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19034_o = n19032_o & n19033_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19035_o = n19031_o | n19034_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19036_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19037_o = n19016_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19038_o = n19036_o & n19037_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19039_o = n19035_o | n19038_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19040_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19041_o = n19016_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19042_o = n19040_o & n19041_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19043_o = n19039_o | n19042_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19044_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19045_o = n19016_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19046_o = n19044_o & n19045_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19047_o = n19043_o | n19046_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19048_o = ~n19047_o;
  /* vlm5030_gl.vhd:2124:34  */
  assign n19050_o = idlat[1];
  /* vlm5030_gl.vhd:2124:25  */
  assign n19051_o = ~n19050_o;
  /* vlm5030_gl.vhd:2124:45  */
  assign n19052_o = idlat[1];
  /* vlm5030_gl.vhd:2124:38  */
  assign n19053_o = {n19051_o, n19052_o};
  /* vlm5030_gl.vhd:2124:60  */
  assign n19054_o = mem1do2ie[2];
  /* vlm5030_gl.vhd:2124:49  */
  assign n19055_o = {n19053_o, n19054_o};
  /* vlm5030_gl.vhd:2124:76  */
  assign n19056_o = mem2do2ie[2];
  /* vlm5030_gl.vhd:2124:65  */
  assign n19057_o = {n19055_o, n19056_o};
  /* vlm5030_gl.vhd:2124:94  */
  assign n19058_o = ieregdrv4ie[2];
  /* vlm5030_gl.vhd:2124:81  */
  assign n19059_o = {n19057_o, n19058_o};
  /* vlm5030_gl.vhd:2124:105  */
  assign n19060_o = i_d[2];
  /* vlm5030_gl.vhd:2124:99  */
  assign n19061_o = {n19059_o, n19060_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19067_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19068_o = n19061_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19069_o = n19067_o & n19068_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19071_o = 1'b0 | n19069_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19073_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19074_o = n19061_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19075_o = n19073_o & n19074_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19076_o = n19071_o | n19075_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19077_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19078_o = n19061_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19079_o = n19077_o & n19078_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19080_o = n19076_o | n19079_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19081_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19082_o = n19061_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19083_o = n19081_o & n19082_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19084_o = n19080_o | n19083_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19085_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19086_o = n19061_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19087_o = n19085_o & n19086_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19088_o = n19084_o | n19087_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19089_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19090_o = n19061_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19091_o = n19089_o & n19090_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19092_o = n19088_o | n19091_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19093_o = ~n19092_o;
  /* vlm5030_gl.vhd:2125:34  */
  assign n19095_o = idlat[2];
  /* vlm5030_gl.vhd:2125:25  */
  assign n19096_o = ~n19095_o;
  /* vlm5030_gl.vhd:2125:45  */
  assign n19097_o = idlat[2];
  /* vlm5030_gl.vhd:2125:38  */
  assign n19098_o = {n19096_o, n19097_o};
  /* vlm5030_gl.vhd:2125:60  */
  assign n19099_o = mem1do2ie[3];
  /* vlm5030_gl.vhd:2125:49  */
  assign n19100_o = {n19098_o, n19099_o};
  /* vlm5030_gl.vhd:2125:76  */
  assign n19101_o = mem2do2ie[3];
  /* vlm5030_gl.vhd:2125:65  */
  assign n19102_o = {n19100_o, n19101_o};
  /* vlm5030_gl.vhd:2125:94  */
  assign n19103_o = ieregdrv4ie[3];
  /* vlm5030_gl.vhd:2125:81  */
  assign n19104_o = {n19102_o, n19103_o};
  /* vlm5030_gl.vhd:2125:105  */
  assign n19105_o = i_d[3];
  /* vlm5030_gl.vhd:2125:99  */
  assign n19106_o = {n19104_o, n19105_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19112_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19113_o = n19106_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19114_o = n19112_o & n19113_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19116_o = 1'b0 | n19114_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19118_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19119_o = n19106_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19120_o = n19118_o & n19119_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19121_o = n19116_o | n19120_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19122_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19123_o = n19106_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19124_o = n19122_o & n19123_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19125_o = n19121_o | n19124_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19126_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19127_o = n19106_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19128_o = n19126_o & n19127_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19129_o = n19125_o | n19128_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19130_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19131_o = n19106_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19132_o = n19130_o & n19131_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19133_o = n19129_o | n19132_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19134_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19135_o = n19106_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19136_o = n19134_o & n19135_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19137_o = n19133_o | n19136_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19138_o = ~n19137_o;
  /* vlm5030_gl.vhd:2126:34  */
  assign n19140_o = idlat[3];
  /* vlm5030_gl.vhd:2126:25  */
  assign n19141_o = ~n19140_o;
  /* vlm5030_gl.vhd:2126:45  */
  assign n19142_o = idlat[3];
  /* vlm5030_gl.vhd:2126:38  */
  assign n19143_o = {n19141_o, n19142_o};
  /* vlm5030_gl.vhd:2126:60  */
  assign n19144_o = mem1do2ie[4];
  /* vlm5030_gl.vhd:2126:49  */
  assign n19145_o = {n19143_o, n19144_o};
  /* vlm5030_gl.vhd:2126:76  */
  assign n19146_o = mem2do2ie[4];
  /* vlm5030_gl.vhd:2126:65  */
  assign n19147_o = {n19145_o, n19146_o};
  /* vlm5030_gl.vhd:2126:94  */
  assign n19148_o = ieregdrv4ie[4];
  /* vlm5030_gl.vhd:2126:81  */
  assign n19149_o = {n19147_o, n19148_o};
  /* vlm5030_gl.vhd:2126:105  */
  assign n19150_o = i_d[4];
  /* vlm5030_gl.vhd:2126:99  */
  assign n19151_o = {n19149_o, n19150_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19157_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19158_o = n19151_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19159_o = n19157_o & n19158_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19161_o = 1'b0 | n19159_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19163_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19164_o = n19151_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19165_o = n19163_o & n19164_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19166_o = n19161_o | n19165_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19167_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19168_o = n19151_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19169_o = n19167_o & n19168_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19170_o = n19166_o | n19169_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19171_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19172_o = n19151_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19173_o = n19171_o & n19172_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19174_o = n19170_o | n19173_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19175_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19176_o = n19151_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19177_o = n19175_o & n19176_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19178_o = n19174_o | n19177_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19179_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19180_o = n19151_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19181_o = n19179_o & n19180_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19182_o = n19178_o | n19181_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19183_o = ~n19182_o;
  /* vlm5030_gl.vhd:2127:34  */
  assign n19185_o = idlat[4];
  /* vlm5030_gl.vhd:2127:25  */
  assign n19186_o = ~n19185_o;
  /* vlm5030_gl.vhd:2127:45  */
  assign n19187_o = idlat[4];
  /* vlm5030_gl.vhd:2127:38  */
  assign n19188_o = {n19186_o, n19187_o};
  /* vlm5030_gl.vhd:2127:60  */
  assign n19189_o = mem1do2ie[5];
  /* vlm5030_gl.vhd:2127:49  */
  assign n19190_o = {n19188_o, n19189_o};
  /* vlm5030_gl.vhd:2127:76  */
  assign n19191_o = mem2do2ie[5];
  /* vlm5030_gl.vhd:2127:65  */
  assign n19192_o = {n19190_o, n19191_o};
  /* vlm5030_gl.vhd:2127:94  */
  assign n19193_o = ieregdrv4ie[5];
  /* vlm5030_gl.vhd:2127:81  */
  assign n19194_o = {n19192_o, n19193_o};
  /* vlm5030_gl.vhd:2127:105  */
  assign n19195_o = i_d[5];
  /* vlm5030_gl.vhd:2127:99  */
  assign n19196_o = {n19194_o, n19195_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19202_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19203_o = n19196_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19204_o = n19202_o & n19203_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19206_o = 1'b0 | n19204_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19208_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19209_o = n19196_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19210_o = n19208_o & n19209_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19211_o = n19206_o | n19210_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19212_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19213_o = n19196_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19214_o = n19212_o & n19213_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19215_o = n19211_o | n19214_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19216_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19217_o = n19196_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19218_o = n19216_o & n19217_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19219_o = n19215_o | n19218_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19220_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19221_o = n19196_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19222_o = n19220_o & n19221_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19223_o = n19219_o | n19222_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19224_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19225_o = n19196_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19226_o = n19224_o & n19225_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19227_o = n19223_o | n19226_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19228_o = ~n19227_o;
  /* vlm5030_gl.vhd:2128:34  */
  assign n19230_o = idlat[5];
  /* vlm5030_gl.vhd:2128:25  */
  assign n19231_o = ~n19230_o;
  /* vlm5030_gl.vhd:2128:45  */
  assign n19232_o = idlat[5];
  /* vlm5030_gl.vhd:2128:38  */
  assign n19233_o = {n19231_o, n19232_o};
  /* vlm5030_gl.vhd:2128:60  */
  assign n19234_o = mem1do2ie[6];
  /* vlm5030_gl.vhd:2128:49  */
  assign n19235_o = {n19233_o, n19234_o};
  /* vlm5030_gl.vhd:2128:76  */
  assign n19236_o = mem2do2ie[6];
  /* vlm5030_gl.vhd:2128:65  */
  assign n19237_o = {n19235_o, n19236_o};
  /* vlm5030_gl.vhd:2128:94  */
  assign n19238_o = ieregdrv4ie[6];
  /* vlm5030_gl.vhd:2128:81  */
  assign n19239_o = {n19237_o, n19238_o};
  /* vlm5030_gl.vhd:2128:105  */
  assign n19240_o = i_d[6];
  /* vlm5030_gl.vhd:2128:99  */
  assign n19241_o = {n19239_o, n19240_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19247_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19248_o = n19241_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19249_o = n19247_o & n19248_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19251_o = 1'b0 | n19249_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19253_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19254_o = n19241_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19255_o = n19253_o & n19254_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19256_o = n19251_o | n19255_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19257_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19258_o = n19241_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19259_o = n19257_o & n19258_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19260_o = n19256_o | n19259_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19261_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19262_o = n19241_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19263_o = n19261_o & n19262_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19264_o = n19260_o | n19263_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19265_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19266_o = n19241_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19267_o = n19265_o & n19266_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19268_o = n19264_o | n19267_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19269_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19270_o = n19241_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19271_o = n19269_o & n19270_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19272_o = n19268_o | n19271_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19273_o = ~n19272_o;
  /* vlm5030_gl.vhd:2129:34  */
  assign n19275_o = idlat[6];
  /* vlm5030_gl.vhd:2129:25  */
  assign n19276_o = ~n19275_o;
  /* vlm5030_gl.vhd:2129:45  */
  assign n19277_o = idlat[6];
  /* vlm5030_gl.vhd:2129:38  */
  assign n19278_o = {n19276_o, n19277_o};
  /* vlm5030_gl.vhd:2129:60  */
  assign n19279_o = mem1do2ie[7];
  /* vlm5030_gl.vhd:2129:49  */
  assign n19280_o = {n19278_o, n19279_o};
  /* vlm5030_gl.vhd:2129:76  */
  assign n19281_o = mem2do2ie[7];
  /* vlm5030_gl.vhd:2129:65  */
  assign n19282_o = {n19280_o, n19281_o};
  /* vlm5030_gl.vhd:2129:94  */
  assign n19283_o = ieregdrv4ie[7];
  /* vlm5030_gl.vhd:2129:81  */
  assign n19284_o = {n19282_o, n19283_o};
  /* vlm5030_gl.vhd:2129:105  */
  assign n19285_o = i_d[7];
  /* vlm5030_gl.vhd:2129:99  */
  assign n19286_o = {n19284_o, n19285_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19292_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19293_o = n19286_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19294_o = n19292_o & n19293_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19296_o = 1'b0 | n19294_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19298_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19299_o = n19286_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19300_o = n19298_o & n19299_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19301_o = n19296_o | n19300_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19302_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19303_o = n19286_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19304_o = n19302_o & n19303_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19305_o = n19301_o | n19304_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19306_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19307_o = n19286_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19308_o = n19306_o & n19307_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19309_o = n19305_o | n19308_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19310_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19311_o = n19286_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19312_o = n19310_o & n19311_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19313_o = n19309_o | n19312_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19314_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19315_o = n19286_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19316_o = n19314_o & n19315_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19317_o = n19313_o | n19316_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19318_o = ~n19317_o;
  /* vlm5030_gl.vhd:2130:34  */
  assign n19320_o = idlat[7];
  /* vlm5030_gl.vhd:2130:25  */
  assign n19321_o = ~n19320_o;
  /* vlm5030_gl.vhd:2130:45  */
  assign n19322_o = idlat[7];
  /* vlm5030_gl.vhd:2130:38  */
  assign n19323_o = {n19321_o, n19322_o};
  /* vlm5030_gl.vhd:2130:60  */
  assign n19324_o = mem1do2ie[8];
  /* vlm5030_gl.vhd:2130:49  */
  assign n19325_o = {n19323_o, n19324_o};
  /* vlm5030_gl.vhd:2130:76  */
  assign n19326_o = mem2do2ie[8];
  /* vlm5030_gl.vhd:2130:65  */
  assign n19327_o = {n19325_o, n19326_o};
  /* vlm5030_gl.vhd:2130:94  */
  assign n19328_o = ieregdrv4ie[8];
  /* vlm5030_gl.vhd:2130:81  */
  assign n19329_o = {n19327_o, n19328_o};
  /* vlm5030_gl.vhd:2130:105  */
  assign n19330_o = i_d[0];
  /* vlm5030_gl.vhd:2130:99  */
  assign n19331_o = {n19329_o, n19330_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19337_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19338_o = n19331_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19339_o = n19337_o & n19338_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19341_o = 1'b0 | n19339_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19343_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19344_o = n19331_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19345_o = n19343_o & n19344_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19346_o = n19341_o | n19345_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19347_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19348_o = n19331_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19349_o = n19347_o & n19348_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19350_o = n19346_o | n19349_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19351_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19352_o = n19331_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19353_o = n19351_o & n19352_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19354_o = n19350_o | n19353_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19355_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19356_o = n19331_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19357_o = n19355_o & n19356_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19358_o = n19354_o | n19357_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19359_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19360_o = n19331_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19361_o = n19359_o & n19360_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19362_o = n19358_o | n19361_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19363_o = ~n19362_o;
  /* vlm5030_gl.vhd:2131:60  */
  assign n19365_o = mem1do2ie[9];
  /* vlm5030_gl.vhd:2131:49  */
  assign n19367_o = {2'b01, n19365_o};
  /* vlm5030_gl.vhd:2131:76  */
  assign n19368_o = mem2do2ie[9];
  /* vlm5030_gl.vhd:2131:65  */
  assign n19369_o = {n19367_o, n19368_o};
  /* vlm5030_gl.vhd:2131:94  */
  assign n19370_o = ieregdrv4ie[9];
  /* vlm5030_gl.vhd:2131:81  */
  assign n19371_o = {n19369_o, n19370_o};
  /* vlm5030_gl.vhd:2131:105  */
  assign n19372_o = i_d[1];
  /* vlm5030_gl.vhd:2131:99  */
  assign n19373_o = {n19371_o, n19372_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19379_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19380_o = n19373_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19381_o = n19379_o & n19380_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19383_o = 1'b0 | n19381_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19385_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19386_o = n19373_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19387_o = n19385_o & n19386_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19388_o = n19383_o | n19387_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19389_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19390_o = n19373_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19391_o = n19389_o & n19390_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19392_o = n19388_o | n19391_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19393_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19394_o = n19373_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19395_o = n19393_o & n19394_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19396_o = n19392_o | n19395_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19397_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19398_o = n19373_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19399_o = n19397_o & n19398_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19400_o = n19396_o | n19399_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19401_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19402_o = n19373_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19403_o = n19401_o & n19402_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19404_o = n19400_o | n19403_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19405_o = ~n19404_o;
  /* vlm5030_gl.vhd:2132:60  */
  assign n19407_o = mem1do2ie[10];
  /* vlm5030_gl.vhd:2132:49  */
  assign n19409_o = {2'b01, n19407_o};
  /* vlm5030_gl.vhd:2132:76  */
  assign n19410_o = mem2do2ie[10];
  /* vlm5030_gl.vhd:2132:65  */
  assign n19411_o = {n19409_o, n19410_o};
  /* vlm5030_gl.vhd:2132:94  */
  assign n19412_o = ieregdrv4ie[10];
  /* vlm5030_gl.vhd:2132:81  */
  assign n19413_o = {n19411_o, n19412_o};
  /* vlm5030_gl.vhd:2132:105  */
  assign n19414_o = i_d[2];
  /* vlm5030_gl.vhd:2132:99  */
  assign n19415_o = {n19413_o, n19414_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19421_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19422_o = n19415_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19423_o = n19421_o & n19422_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19425_o = 1'b0 | n19423_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19427_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19428_o = n19415_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19429_o = n19427_o & n19428_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19430_o = n19425_o | n19429_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19431_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19432_o = n19415_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19433_o = n19431_o & n19432_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19434_o = n19430_o | n19433_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19435_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19436_o = n19415_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19437_o = n19435_o & n19436_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19438_o = n19434_o | n19437_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19439_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19440_o = n19415_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19441_o = n19439_o & n19440_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19442_o = n19438_o | n19441_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19443_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19444_o = n19415_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19445_o = n19443_o & n19444_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19446_o = n19442_o | n19445_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19447_o = ~n19446_o;
  /* vlm5030_gl.vhd:2133:60  */
  assign n19449_o = mem1do2ie[11];
  /* vlm5030_gl.vhd:2133:49  */
  assign n19451_o = {2'b01, n19449_o};
  /* vlm5030_gl.vhd:2133:76  */
  assign n19452_o = mem2do2ie[11];
  /* vlm5030_gl.vhd:2133:65  */
  assign n19453_o = {n19451_o, n19452_o};
  /* vlm5030_gl.vhd:2133:94  */
  assign n19454_o = ieregdrv4ie[11];
  /* vlm5030_gl.vhd:2133:81  */
  assign n19455_o = {n19453_o, n19454_o};
  /* vlm5030_gl.vhd:2133:105  */
  assign n19456_o = i_d[3];
  /* vlm5030_gl.vhd:2133:99  */
  assign n19457_o = {n19455_o, n19456_o};
  /* vlm5030_pack.vhd:50:26  */
  assign n19463_o = nie_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19464_o = n19457_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19465_o = n19463_o & n19464_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19467_o = 1'b0 | n19465_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19469_o = nie_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19470_o = n19457_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19471_o = n19469_o & n19470_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19472_o = n19467_o | n19471_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19473_o = nie_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19474_o = n19457_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19475_o = n19473_o & n19474_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19476_o = n19472_o | n19475_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19477_o = nie_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19478_o = n19457_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19479_o = n19477_o & n19478_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19480_o = n19476_o | n19479_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19481_o = nie_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19482_o = n19457_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19483_o = n19481_o & n19482_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19484_o = n19480_o | n19483_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19485_o = nie_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19486_o = n19457_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19487_o = n19485_o & n19486_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19488_o = n19484_o | n19487_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19489_o = ~n19488_o;
  /* vlm5030_gl.vhd:2143:12  */
  assign dac_block_pwmsel = n19592_o; // (signal)
  /* vlm5030_gl.vhd:2147:14  */
  assign dac_block_pwm_block_pwm0 = n19500_o; // (signal)
  /* vlm5030_gl.vhd:2147:20  */
  assign dac_block_pwm_block_pwm1 = n19496_o; // (signal)
  /* vlm5030_gl.vhd:2147:26  */
  assign dac_block_pwm_block_pwm2 = n19492_o; // (signal)
  /* vlm5030_gl.vhd:2149:14  */
  assign dac_block_pwm_block_nc2d10xr9del = dac_block_pwm_block_nc2d10xr9del_b_o_out; // (signal)
  /* vlm5030_gl.vhd:2153:14  */
  assign dac_block_pwm_block_pwmreg1toggle = dac_block_pwm_block_pwmreg0; // (signal)
  /* vlm5030_gl.vhd:2154:14  */
  assign dac_block_pwm_block_pwmreg2toggle = n19510_o; // (signal)
  /* vlm5030_gl.vhd:2155:14  */
  assign dac_block_pwm_block_pwmreg0 = n19595_q; // (signal)
  /* vlm5030_gl.vhd:2155:23  */
  assign dac_block_pwm_block_pwmreg1 = n19597_q; // (signal)
  /* vlm5030_gl.vhd:2156:14  */
  assign dac_block_pwm_block_pwmreg2 = n19599_q; // (signal)
  /* vlm5030_gl.vhd:2158:14  */
  assign dac_block_pwm_block_pwmcomm = n19554_o; // (signal)
  /* vlm5030_gl.vhd:2159:14  */
  assign dac_block_pwm_block_pwmcommdel = dac_block_pwm_block_pwmcommdel_b_o_out; // (signal)
  /* vlm5030_gl.vhd:2160:14  */
  assign dac_block_pwm_block_pwmcommand = n19560_o; // (signal)
  /* vlm5030_gl.vhd:2161:14  */
  assign dac_block_pwm_block_pwmcomp = n19588_o; // (signal)
  /* vlm5030_gl.vhd:2165:24  */
  assign n19490_o = ieaddrreg[4];
  /* vlm5030_gl.vhd:2165:45  */
  assign n19491_o = ~tstenie2dac;
  /* vlm5030_gl.vhd:2165:28  */
  assign n19492_o = n19491_o ? n19490_o : n19493_o;
  /* vlm5030_gl.vhd:2165:59  */
  assign n19493_o = nie[4];
  /* vlm5030_gl.vhd:2166:24  */
  assign n19494_o = ieaddrreg[3];
  /* vlm5030_gl.vhd:2166:45  */
  assign n19495_o = ~tstenie2dac;
  /* vlm5030_gl.vhd:2166:28  */
  assign n19496_o = n19495_o ? n19494_o : n19497_o;
  /* vlm5030_gl.vhd:2166:59  */
  assign n19497_o = nie[3];
  /* vlm5030_gl.vhd:2167:24  */
  assign n19498_o = ieaddrreg[2];
  /* vlm5030_gl.vhd:2167:45  */
  assign n19499_o = ~tstenie2dac;
  /* vlm5030_gl.vhd:2167:28  */
  assign n19500_o = n19499_o ? n19498_o : n19501_o;
  /* vlm5030_gl.vhd:2167:59  */
  assign n19501_o = nie[2];
  /* vlm5030_gl.vhd:2169:7  */
  vlm5030_delay_inv_4 dac_block_pwm_block_nc2d10xr9del_b (
    .i_clk_base(n19502_o),
    .i_clk_val(n19503_o),
    .i_clk_rise(n19504_o),
    .i_clk_fall(n19505_o),
    .i_in(n19506_o),
    .o_out(dac_block_pwm_block_nc2d10xr9del_b_o_out));
  assign n19502_o = osc[0];
  assign n19503_o = osc[1];
  assign n19504_o = osc[2];
  assign n19505_o = osc[3];
  /* vlm5030_gl.vhd:2176:29  */
  assign n19506_o = c2d10xr9[1];
  /* vlm5030_gl.vhd:2183:25  */
  assign n19508_o = ~dac_block_pwm_block_pwmreg1;
  /* vlm5030_gl.vhd:2183:43  */
  assign n19509_o = ~dac_block_pwm_block_pwmreg0;
  /* vlm5030_gl.vhd:2183:38  */
  assign n19510_o = ~(n19508_o | n19509_o);
  assign n19518_o = clk2gd5[0];
  /* clock_functions_pack.vhd:65:42  */
  assign n19520_o = clk2gd5[2];
  /* vlm5030_gl.vhd:2188:27  */
  assign n19522_o = ~dac_block_pwm_block_nc2d10xr9del;
  /* vlm5030_gl.vhd:2195:24  */
  assign n19523_o = ~dac_block_pwm_block_pwmreg0;
  /* vlm5030_gl.vhd:2197:26  */
  assign n19524_o = ~dac_block_pwm_block_pwmreg1;
  /* vlm5030_gl.vhd:2196:13  */
  assign n19525_o = dac_block_pwm_block_pwmreg1toggle ? n19524_o : dac_block_pwm_block_pwmreg1;
  /* vlm5030_gl.vhd:2200:26  */
  assign n19526_o = ~dac_block_pwm_block_pwmreg2;
  /* vlm5030_gl.vhd:2199:13  */
  assign n19527_o = dac_block_pwm_block_pwmreg2toggle ? n19526_o : dac_block_pwm_block_pwmreg2;
  /* vlm5030_gl.vhd:2188:11  */
  assign n19529_o = n19522_o ? 1'b0 : n19523_o;
  /* vlm5030_gl.vhd:2188:11  */
  assign n19531_o = n19522_o ? 1'b0 : n19525_o;
  /* vlm5030_gl.vhd:2188:11  */
  assign n19533_o = n19522_o ? 1'b0 : n19527_o;
  /* vlm5030_gl.vhd:2207:31  */
  assign n19539_o = {dac_block_pwm_block_pwmreg0, dac_block_pwm_block_pwmreg1};
  /* vlm5030_gl.vhd:2207:41  */
  assign n19540_o = {n19539_o, dac_block_pwm_block_pwmreg2};
  /* vlm5030_pack.vhd:40:24  */
  assign n19546_o = n19540_o[2];
  /* vlm5030_pack.vhd:40:20  */
  assign n19548_o = 1'b0 | n19546_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n19550_o = n19540_o[1];
  /* vlm5030_pack.vhd:40:20  */
  assign n19551_o = n19548_o | n19550_o;
  /* vlm5030_pack.vhd:40:24  */
  assign n19552_o = n19540_o[0];
  /* vlm5030_pack.vhd:40:20  */
  assign n19553_o = n19551_o | n19552_o;
  /* vlm5030_pack.vhd:42:12  */
  assign n19554_o = ~n19553_o;
  /* vlm5030_gl.vhd:2208:7  */
  vlm5030_delay_4 dac_block_pwm_block_pwmcommdel_b (
    .i_clk_base(n19555_o),
    .i_clk_val(n19556_o),
    .i_clk_rise(n19557_o),
    .i_clk_fall(n19558_o),
    .i_in(dac_block_pwm_block_pwmcomm),
    .o_out(dac_block_pwm_block_pwmcommdel_b_o_out));
  assign n19555_o = osc[0];
  assign n19556_o = osc[1];
  assign n19557_o = osc[2];
  assign n19558_o = osc[3];
  /* vlm5030_gl.vhd:2218:29  */
  assign n19560_o = dac_block_pwm_block_pwmcomm & dac_block_pwm_block_pwmcommdel;
  /* vlm5030_gl.vhd:2220:29  */
  assign n19562_o = {dac_block_pwm_block_pwm2, dac_block_pwm_block_pwm1};
  /* vlm5030_gl.vhd:2220:36  */
  assign n19563_o = {n19562_o, dac_block_pwm_block_pwm0};
  /* vlm5030_gl.vhd:2220:52  */
  assign n19564_o = {dac_block_pwm_block_pwmreg2, dac_block_pwm_block_pwmreg1};
  /* vlm5030_gl.vhd:2220:62  */
  assign n19565_o = {n19564_o, dac_block_pwm_block_pwmreg0};
  /* vlm5030_pack.vhd:60:26  */
  assign n19571_o = n19563_o[2];
  /* vlm5030_pack.vhd:60:43  */
  assign n19572_o = n19565_o[2];
  /* vlm5030_pack.vhd:60:36  */
  assign n19573_o = ~n19572_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n19574_o = n19571_o & n19573_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n19576_o = 1'b0 | n19574_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n19578_o = n19563_o[1];
  /* vlm5030_pack.vhd:60:43  */
  assign n19579_o = n19565_o[1];
  /* vlm5030_pack.vhd:60:36  */
  assign n19580_o = ~n19579_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n19581_o = n19578_o & n19580_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n19582_o = n19576_o | n19581_o;
  /* vlm5030_pack.vhd:60:26  */
  assign n19583_o = n19563_o[0];
  /* vlm5030_pack.vhd:60:43  */
  assign n19584_o = n19565_o[0];
  /* vlm5030_pack.vhd:60:36  */
  assign n19585_o = ~n19584_o;
  /* vlm5030_pack.vhd:60:32  */
  assign n19586_o = n19583_o & n19585_o;
  /* vlm5030_pack.vhd:60:20  */
  assign n19587_o = n19582_o | n19586_o;
  /* vlm5030_pack.vhd:62:12  */
  assign n19588_o = ~n19587_o;
  /* vlm5030_gl.vhd:2222:7  */
  vlm5030_srlatch dac_block_pwm_block_pwmsr_b (
    .i_clk(n19589_o),
    .i_res(dac_block_pwm_block_pwmcomp),
    .i_set(dac_block_pwm_block_pwmcommand),
    .o_q(dac_block_pwm_block_pwmsr_b_o_q));
  /* vlm5030_gl.vhd:2224:24  */
  assign n19589_o = osc[0];
  /* vlm5030_gl.vhd:2229:17  */
  assign n19591_o = ~i_vcu;
  /* vlm5030_gl.vhd:2229:27  */
  assign n19592_o = tstenie2dac ? n19591_o : n19593_o;
  /* vlm5030_gl.vhd:2230:17  */
  assign n19593_o = ~pwmsr;
  /* vlm5030_gl.vhd:2187:9  */
  assign n19594_o = n19520_o ? n19529_o : dac_block_pwm_block_pwmreg0;
  /* vlm5030_gl.vhd:2187:9  */
  always @(posedge n19518_o)
    n19595_q <= n19594_o;
  /* vlm5030_gl.vhd:2187:9  */
  assign n19596_o = n19520_o ? n19531_o : dac_block_pwm_block_pwmreg1;
  /* vlm5030_gl.vhd:2187:9  */
  always @(posedge n19518_o)
    n19597_q <= n19596_o;
  /* vlm5030_gl.vhd:2187:9  */
  assign n19598_o = n19520_o ? n19533_o : dac_block_pwm_block_pwmreg2;
  /* vlm5030_gl.vhd:2187:9  */
  always @(posedge n19518_o)
    n19599_q <= n19598_o;
  /* vlm5030_gl.vhd:2235:14  */
  assign dac_block_dacrom_block_ndac = n19605_o; // (signal)
  /* vlm5030_gl.vhd:2236:14  */
  assign dac_block_dacrom_block_dacval = n19615_o; // (signal)
  /* vlm5030_gl.vhd:2236:22  */
  assign dac_block_dacrom_block_dacpwm = n19616_o; // (signal)
  /* vlm5030_gl.vhd:2239:24  */
  assign n19600_o = ieaddrreg[9];
  /* vlm5030_gl.vhd:2239:43  */
  assign n19601_o = ieaddrreg[8:5];
  /* vlm5030_gl.vhd:2239:30  */
  assign n19602_o = ~n19601_o;
  /* vlm5030_gl.vhd:2239:28  */
  assign n19603_o = {n19600_o, n19602_o};
  /* vlm5030_gl.vhd:2239:73  */
  assign n19604_o = ~tstenie2dac;
  /* vlm5030_gl.vhd:2239:56  */
  assign n19605_o = n19604_o ? n19603_o : n19609_o;
  /* vlm5030_gl.vhd:2240:18  */
  assign n19606_o = nie[9];
  /* vlm5030_gl.vhd:2240:31  */
  assign n19607_o = nie[8:5];
  /* vlm5030_gl.vhd:2240:24  */
  assign n19608_o = ~n19607_o;
  /* vlm5030_gl.vhd:2240:22  */
  assign n19609_o = {n19606_o, n19608_o};
  /* vlm5030_gl.vhd:2248:31  */
  assign n19610_o = ~dac_block_dacrom_block_ndac;
  /* vlm5030_gl.vhd:2248:17  */
  assign n19611_o = {{2{n19610_o[4]}}, n19610_o}; // sext
  /* vlm5030_gl.vhd:2248:57  */
  assign n19613_o = n19611_o + 7'b0010000;
  /* vlm5030_gl.vhd:2248:61  */
  assign n19615_o = n19613_o + 7'b0000001;
  /* vlm5030_gl.vhd:2250:24  */
  assign n19616_o = dac_block_pwmsel ? dac_block_dacrom_block_dacval : n19618_o;
  /* vlm5030_gl.vhd:2250:54  */
  assign n19618_o = dac_block_dacrom_block_dacval + 7'b0000001;
  /* vlm5030_gl.vhd:2252:39  */
  assign n19619_o = dac_block_dacrom_block_dacpwm[5:0];
  /* vlm5030_gl.vhd:2266:12  */
  assign abus_block_wl = n19625_o; // (signal)
  /* vlm5030_gl.vhd:2269:36  */
  assign n19621_o = {eaoen, enie2a};
  /* vlm5030_gl.vhd:2269:55  */
  assign n19622_o = {n19621_o, tstenid2a};
  /* vlm5030_gl.vhd:2269:68  */
  assign n19623_o = {n19622_o, tstenie2a};
  /* vlm5030_gl.vhd:2269:82  */
  assign n19624_o = {n19623_o, tstenctrl2a};
  /* vlm5030_gl.vhd:2269:96  */
  assign n19625_o = {n19624_o, tstenie2dac};
  /* vlm5030_gl.vhd:2271:31  */
  assign n19627_o = aq[0];
  /* vlm5030_gl.vhd:2271:49  */
  assign n19628_o = ieaddrreg[0];
  /* vlm5030_gl.vhd:2271:36  */
  assign n19629_o = {n19627_o, n19628_o};
  /* vlm5030_gl.vhd:2271:64  */
  assign n19630_o = nid[0];
  /* vlm5030_gl.vhd:2271:57  */
  assign n19631_o = ~n19630_o;
  /* vlm5030_gl.vhd:2271:55  */
  assign n19632_o = {n19629_o, n19631_o};
  /* vlm5030_gl.vhd:2271:77  */
  assign n19633_o = nie[0];
  /* vlm5030_gl.vhd:2271:70  */
  assign n19634_o = ~n19633_o;
  /* vlm5030_gl.vhd:2271:68  */
  assign n19635_o = {n19632_o, n19634_o};
  /* vlm5030_gl.vhd:2271:82  */
  assign n19637_o = {n19635_o, 1'b0};
  /* vlm5030_gl.vhd:2271:96  */
  assign n19639_o = {n19637_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n19645_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19646_o = n19639_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19647_o = n19645_o & n19646_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19649_o = 1'b0 | n19647_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19651_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19652_o = n19639_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19653_o = n19651_o & n19652_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19654_o = n19649_o | n19653_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19655_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19656_o = n19639_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19657_o = n19655_o & n19656_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19658_o = n19654_o | n19657_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19659_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19660_o = n19639_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19661_o = n19659_o & n19660_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19662_o = n19658_o | n19661_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19663_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19664_o = n19639_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19665_o = n19663_o & n19664_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19666_o = n19662_o | n19665_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19667_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19668_o = n19639_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19669_o = n19667_o & n19668_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19670_o = n19666_o | n19669_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19671_o = ~n19670_o;
  /* vlm5030_gl.vhd:2271:16  */
  assign n19672_o = ~n19671_o;
  /* vlm5030_gl.vhd:2272:31  */
  assign n19674_o = aq[1];
  /* vlm5030_gl.vhd:2272:49  */
  assign n19675_o = ieaddrreg[1];
  /* vlm5030_gl.vhd:2272:36  */
  assign n19676_o = {n19674_o, n19675_o};
  /* vlm5030_gl.vhd:2272:64  */
  assign n19677_o = nid[1];
  /* vlm5030_gl.vhd:2272:57  */
  assign n19678_o = ~n19677_o;
  /* vlm5030_gl.vhd:2272:55  */
  assign n19679_o = {n19676_o, n19678_o};
  /* vlm5030_gl.vhd:2272:77  */
  assign n19680_o = nie[1];
  /* vlm5030_gl.vhd:2272:70  */
  assign n19681_o = ~n19680_o;
  /* vlm5030_gl.vhd:2272:68  */
  assign n19682_o = {n19679_o, n19681_o};
  /* vlm5030_gl.vhd:2272:82  */
  assign n19684_o = {n19682_o, 1'b0};
  /* vlm5030_gl.vhd:2272:96  */
  assign n19686_o = {n19684_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n19692_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19693_o = n19686_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19694_o = n19692_o & n19693_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19696_o = 1'b0 | n19694_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19698_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19699_o = n19686_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19700_o = n19698_o & n19699_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19701_o = n19696_o | n19700_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19702_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19703_o = n19686_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19704_o = n19702_o & n19703_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19705_o = n19701_o | n19704_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19706_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19707_o = n19686_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19708_o = n19706_o & n19707_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19709_o = n19705_o | n19708_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19710_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19711_o = n19686_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19712_o = n19710_o & n19711_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19713_o = n19709_o | n19712_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19714_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19715_o = n19686_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19716_o = n19714_o & n19715_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19717_o = n19713_o | n19716_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19718_o = ~n19717_o;
  /* vlm5030_gl.vhd:2272:16  */
  assign n19719_o = ~n19718_o;
  /* vlm5030_gl.vhd:2273:31  */
  assign n19721_o = aq[2];
  /* vlm5030_gl.vhd:2273:49  */
  assign n19722_o = ieaddrreg[2];
  /* vlm5030_gl.vhd:2273:36  */
  assign n19723_o = {n19721_o, n19722_o};
  /* vlm5030_gl.vhd:2273:64  */
  assign n19724_o = nid[2];
  /* vlm5030_gl.vhd:2273:57  */
  assign n19725_o = ~n19724_o;
  /* vlm5030_gl.vhd:2273:55  */
  assign n19726_o = {n19723_o, n19725_o};
  /* vlm5030_gl.vhd:2273:77  */
  assign n19727_o = nie[2];
  /* vlm5030_gl.vhd:2273:70  */
  assign n19728_o = ~n19727_o;
  /* vlm5030_gl.vhd:2273:68  */
  assign n19729_o = {n19726_o, n19728_o};
  /* vlm5030_gl.vhd:2273:82  */
  assign n19731_o = {n19729_o, 1'b0};
  /* vlm5030_gl.vhd:2273:96  */
  assign n19733_o = {n19731_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n19739_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19740_o = n19733_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19741_o = n19739_o & n19740_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19743_o = 1'b0 | n19741_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19745_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19746_o = n19733_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19747_o = n19745_o & n19746_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19748_o = n19743_o | n19747_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19749_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19750_o = n19733_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19751_o = n19749_o & n19750_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19752_o = n19748_o | n19751_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19753_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19754_o = n19733_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19755_o = n19753_o & n19754_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19756_o = n19752_o | n19755_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19757_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19758_o = n19733_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19759_o = n19757_o & n19758_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19760_o = n19756_o | n19759_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19761_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19762_o = n19733_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19763_o = n19761_o & n19762_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19764_o = n19760_o | n19763_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19765_o = ~n19764_o;
  /* vlm5030_gl.vhd:2273:16  */
  assign n19766_o = ~n19765_o;
  /* vlm5030_gl.vhd:2274:31  */
  assign n19768_o = aq[3];
  /* vlm5030_gl.vhd:2274:49  */
  assign n19769_o = ieaddrreg[3];
  /* vlm5030_gl.vhd:2274:36  */
  assign n19770_o = {n19768_o, n19769_o};
  /* vlm5030_gl.vhd:2274:64  */
  assign n19771_o = nid[3];
  /* vlm5030_gl.vhd:2274:57  */
  assign n19772_o = ~n19771_o;
  /* vlm5030_gl.vhd:2274:55  */
  assign n19773_o = {n19770_o, n19772_o};
  /* vlm5030_gl.vhd:2274:77  */
  assign n19774_o = nie[3];
  /* vlm5030_gl.vhd:2274:70  */
  assign n19775_o = ~n19774_o;
  /* vlm5030_gl.vhd:2274:68  */
  assign n19776_o = {n19773_o, n19775_o};
  /* vlm5030_gl.vhd:2274:82  */
  assign n19778_o = {n19776_o, 1'b0};
  /* vlm5030_gl.vhd:2274:96  */
  assign n19780_o = {n19778_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n19786_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19787_o = n19780_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19788_o = n19786_o & n19787_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19790_o = 1'b0 | n19788_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19792_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19793_o = n19780_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19794_o = n19792_o & n19793_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19795_o = n19790_o | n19794_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19796_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19797_o = n19780_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19798_o = n19796_o & n19797_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19799_o = n19795_o | n19798_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19800_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19801_o = n19780_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19802_o = n19800_o & n19801_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19803_o = n19799_o | n19802_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19804_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19805_o = n19780_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19806_o = n19804_o & n19805_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19807_o = n19803_o | n19806_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19808_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19809_o = n19780_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19810_o = n19808_o & n19809_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19811_o = n19807_o | n19810_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19812_o = ~n19811_o;
  /* vlm5030_gl.vhd:2274:16  */
  assign n19813_o = ~n19812_o;
  /* vlm5030_gl.vhd:2275:31  */
  assign n19815_o = aq[4];
  /* vlm5030_gl.vhd:2275:49  */
  assign n19816_o = ieaddrreg[4];
  /* vlm5030_gl.vhd:2275:36  */
  assign n19817_o = {n19815_o, n19816_o};
  /* vlm5030_gl.vhd:2275:64  */
  assign n19818_o = nid[4];
  /* vlm5030_gl.vhd:2275:57  */
  assign n19819_o = ~n19818_o;
  /* vlm5030_gl.vhd:2275:55  */
  assign n19820_o = {n19817_o, n19819_o};
  /* vlm5030_gl.vhd:2275:77  */
  assign n19821_o = nie[4];
  /* vlm5030_gl.vhd:2275:70  */
  assign n19822_o = ~n19821_o;
  /* vlm5030_gl.vhd:2275:68  */
  assign n19823_o = {n19820_o, n19822_o};
  /* vlm5030_gl.vhd:2275:82  */
  assign n19825_o = {n19823_o, 1'b0};
  /* vlm5030_gl.vhd:2275:96  */
  assign n19827_o = {n19825_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n19833_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19834_o = n19827_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19835_o = n19833_o & n19834_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19837_o = 1'b0 | n19835_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19839_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19840_o = n19827_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19841_o = n19839_o & n19840_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19842_o = n19837_o | n19841_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19843_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19844_o = n19827_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19845_o = n19843_o & n19844_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19846_o = n19842_o | n19845_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19847_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19848_o = n19827_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19849_o = n19847_o & n19848_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19850_o = n19846_o | n19849_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19851_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19852_o = n19827_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19853_o = n19851_o & n19852_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19854_o = n19850_o | n19853_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19855_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19856_o = n19827_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19857_o = n19855_o & n19856_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19858_o = n19854_o | n19857_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19859_o = ~n19858_o;
  /* vlm5030_gl.vhd:2275:16  */
  assign n19860_o = ~n19859_o;
  /* vlm5030_gl.vhd:2276:31  */
  assign n19862_o = aq[5];
  /* vlm5030_gl.vhd:2276:49  */
  assign n19863_o = ieaddrreg[5];
  /* vlm5030_gl.vhd:2276:36  */
  assign n19864_o = {n19862_o, n19863_o};
  /* vlm5030_gl.vhd:2276:64  */
  assign n19865_o = nid[5];
  /* vlm5030_gl.vhd:2276:57  */
  assign n19866_o = ~n19865_o;
  /* vlm5030_gl.vhd:2276:55  */
  assign n19867_o = {n19864_o, n19866_o};
  /* vlm5030_gl.vhd:2276:77  */
  assign n19868_o = nie[5];
  /* vlm5030_gl.vhd:2276:70  */
  assign n19869_o = ~n19868_o;
  /* vlm5030_gl.vhd:2276:68  */
  assign n19870_o = {n19867_o, n19869_o};
  /* vlm5030_gl.vhd:2276:82  */
  assign n19872_o = {n19870_o, 1'b0};
  /* vlm5030_gl.vhd:2276:96  */
  assign n19874_o = {n19872_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n19880_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19881_o = n19874_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19882_o = n19880_o & n19881_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19884_o = 1'b0 | n19882_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19886_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19887_o = n19874_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19888_o = n19886_o & n19887_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19889_o = n19884_o | n19888_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19890_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19891_o = n19874_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19892_o = n19890_o & n19891_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19893_o = n19889_o | n19892_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19894_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19895_o = n19874_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19896_o = n19894_o & n19895_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19897_o = n19893_o | n19896_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19898_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19899_o = n19874_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19900_o = n19898_o & n19899_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19901_o = n19897_o | n19900_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19902_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19903_o = n19874_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19904_o = n19902_o & n19903_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19905_o = n19901_o | n19904_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19906_o = ~n19905_o;
  /* vlm5030_gl.vhd:2276:16  */
  assign n19907_o = ~n19906_o;
  /* vlm5030_gl.vhd:2277:31  */
  assign n19909_o = aq[6];
  /* vlm5030_gl.vhd:2277:49  */
  assign n19910_o = ieaddrreg[6];
  /* vlm5030_gl.vhd:2277:36  */
  assign n19911_o = {n19909_o, n19910_o};
  /* vlm5030_gl.vhd:2277:64  */
  assign n19912_o = nid[6];
  /* vlm5030_gl.vhd:2277:57  */
  assign n19913_o = ~n19912_o;
  /* vlm5030_gl.vhd:2277:55  */
  assign n19914_o = {n19911_o, n19913_o};
  /* vlm5030_gl.vhd:2277:77  */
  assign n19915_o = nie[6];
  /* vlm5030_gl.vhd:2277:70  */
  assign n19916_o = ~n19915_o;
  /* vlm5030_gl.vhd:2277:68  */
  assign n19917_o = {n19914_o, n19916_o};
  /* vlm5030_gl.vhd:2277:82  */
  assign n19919_o = {n19917_o, 1'b0};
  /* vlm5030_gl.vhd:2277:96  */
  assign n19921_o = {n19919_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n19927_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19928_o = n19921_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19929_o = n19927_o & n19928_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19931_o = 1'b0 | n19929_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19933_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19934_o = n19921_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19935_o = n19933_o & n19934_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19936_o = n19931_o | n19935_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19937_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19938_o = n19921_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19939_o = n19937_o & n19938_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19940_o = n19936_o | n19939_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19941_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19942_o = n19921_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19943_o = n19941_o & n19942_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19944_o = n19940_o | n19943_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19945_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19946_o = n19921_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19947_o = n19945_o & n19946_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19948_o = n19944_o | n19947_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19949_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19950_o = n19921_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19951_o = n19949_o & n19950_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19952_o = n19948_o | n19951_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n19953_o = ~n19952_o;
  /* vlm5030_gl.vhd:2277:16  */
  assign n19954_o = ~n19953_o;
  /* vlm5030_gl.vhd:2278:31  */
  assign n19956_o = aq[7];
  /* vlm5030_gl.vhd:2278:49  */
  assign n19957_o = ieaddrreg[7];
  /* vlm5030_gl.vhd:2278:36  */
  assign n19958_o = {n19956_o, n19957_o};
  /* vlm5030_gl.vhd:2278:64  */
  assign n19959_o = nid[7];
  /* vlm5030_gl.vhd:2278:57  */
  assign n19960_o = ~n19959_o;
  /* vlm5030_gl.vhd:2278:55  */
  assign n19961_o = {n19958_o, n19960_o};
  /* vlm5030_gl.vhd:2278:77  */
  assign n19962_o = nie[7];
  /* vlm5030_gl.vhd:2278:70  */
  assign n19963_o = ~n19962_o;
  /* vlm5030_gl.vhd:2278:68  */
  assign n19964_o = {n19961_o, n19963_o};
  /* vlm5030_gl.vhd:2278:82  */
  assign n19966_o = {n19964_o, 1'b0};
  /* vlm5030_gl.vhd:2278:96  */
  assign n19968_o = {n19966_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n19974_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n19975_o = n19968_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n19976_o = n19974_o & n19975_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19978_o = 1'b0 | n19976_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19980_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n19981_o = n19968_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n19982_o = n19980_o & n19981_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19983_o = n19978_o | n19982_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19984_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n19985_o = n19968_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n19986_o = n19984_o & n19985_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19987_o = n19983_o | n19986_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19988_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n19989_o = n19968_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n19990_o = n19988_o & n19989_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19991_o = n19987_o | n19990_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19992_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n19993_o = n19968_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n19994_o = n19992_o & n19993_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19995_o = n19991_o | n19994_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n19996_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n19997_o = n19968_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n19998_o = n19996_o & n19997_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n19999_o = n19995_o | n19998_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20000_o = ~n19999_o;
  /* vlm5030_gl.vhd:2278:16  */
  assign n20001_o = ~n20000_o;
  /* vlm5030_gl.vhd:2279:31  */
  assign n20003_o = aq[8];
  /* vlm5030_gl.vhd:2279:49  */
  assign n20004_o = ieaddrreg[8];
  /* vlm5030_gl.vhd:2279:36  */
  assign n20005_o = {n20003_o, n20004_o};
  /* vlm5030_gl.vhd:2279:64  */
  assign n20006_o = nid[8];
  /* vlm5030_gl.vhd:2279:57  */
  assign n20007_o = ~n20006_o;
  /* vlm5030_gl.vhd:2279:55  */
  assign n20008_o = {n20005_o, n20007_o};
  /* vlm5030_gl.vhd:2279:77  */
  assign n20009_o = nie[8];
  /* vlm5030_gl.vhd:2279:70  */
  assign n20010_o = ~n20009_o;
  /* vlm5030_gl.vhd:2279:68  */
  assign n20011_o = {n20008_o, n20010_o};
  /* vlm5030_gl.vhd:2279:82  */
  assign n20013_o = {n20011_o, 1'b0};
  /* vlm5030_gl.vhd:2279:96  */
  assign n20015_o = {n20013_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n20021_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n20022_o = n20015_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n20023_o = n20021_o & n20022_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20025_o = 1'b0 | n20023_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20027_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n20028_o = n20015_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n20029_o = n20027_o & n20028_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20030_o = n20025_o | n20029_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20031_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n20032_o = n20015_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n20033_o = n20031_o & n20032_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20034_o = n20030_o | n20033_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20035_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n20036_o = n20015_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n20037_o = n20035_o & n20036_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20038_o = n20034_o | n20037_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20039_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n20040_o = n20015_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n20041_o = n20039_o & n20040_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20042_o = n20038_o | n20041_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20043_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n20044_o = n20015_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n20045_o = n20043_o & n20044_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20046_o = n20042_o | n20045_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20047_o = ~n20046_o;
  /* vlm5030_gl.vhd:2279:16  */
  assign n20048_o = ~n20047_o;
  /* vlm5030_gl.vhd:2280:31  */
  assign n20050_o = aq[9];
  /* vlm5030_gl.vhd:2280:51  */
  assign n20051_o = ieaddrreg[9];
  /* vlm5030_gl.vhd:2280:38  */
  assign n20052_o = ~n20051_o;
  /* vlm5030_gl.vhd:2280:36  */
  assign n20053_o = {n20050_o, n20052_o};
  /* vlm5030_gl.vhd:2280:64  */
  assign n20054_o = nid[9];
  /* vlm5030_gl.vhd:2280:57  */
  assign n20055_o = ~n20054_o;
  /* vlm5030_gl.vhd:2280:55  */
  assign n20056_o = {n20053_o, n20055_o};
  /* vlm5030_gl.vhd:2280:77  */
  assign n20057_o = nie[9];
  /* vlm5030_gl.vhd:2280:70  */
  assign n20058_o = ~n20057_o;
  /* vlm5030_gl.vhd:2280:68  */
  assign n20059_o = {n20056_o, n20058_o};
  /* vlm5030_gl.vhd:2280:82  */
  assign n20061_o = {n20059_o, 1'b0};
  /* vlm5030_gl.vhd:2280:96  */
  assign n20063_o = {n20061_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n20069_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n20070_o = n20063_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n20071_o = n20069_o & n20070_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20073_o = 1'b0 | n20071_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20075_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n20076_o = n20063_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n20077_o = n20075_o & n20076_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20078_o = n20073_o | n20077_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20079_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n20080_o = n20063_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n20081_o = n20079_o & n20080_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20082_o = n20078_o | n20081_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20083_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n20084_o = n20063_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n20085_o = n20083_o & n20084_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20086_o = n20082_o | n20085_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20087_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n20088_o = n20063_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n20089_o = n20087_o & n20088_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20090_o = n20086_o | n20089_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20091_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n20092_o = n20063_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n20093_o = n20091_o & n20092_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20094_o = n20090_o | n20093_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20095_o = ~n20094_o;
  /* vlm5030_gl.vhd:2280:16  */
  assign n20096_o = ~n20095_o;
  /* vlm5030_gl.vhd:2281:31  */
  assign n20098_o = aq[10];
  /* vlm5030_gl.vhd:2281:36  */
  assign n20099_o = {n20098_o, pitchoverflow};
  /* vlm5030_gl.vhd:2281:55  */
  assign n20101_o = {n20099_o, 1'b0};
  /* vlm5030_gl.vhd:2281:68  */
  assign n20103_o = {n20101_o, 1'b0};
  /* vlm5030_gl.vhd:2281:90  */
  assign n20104_o = c2d0[1];
  /* vlm5030_gl.vhd:2281:82  */
  assign n20105_o = {n20103_o, n20104_o};
  /* vlm5030_gl.vhd:2281:96  */
  assign n20106_o = {n20105_o, pwmsr};
  /* vlm5030_pack.vhd:50:26  */
  assign n20112_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n20113_o = n20106_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n20114_o = n20112_o & n20113_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20116_o = 1'b0 | n20114_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20118_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n20119_o = n20106_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n20120_o = n20118_o & n20119_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20121_o = n20116_o | n20120_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20122_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n20123_o = n20106_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n20124_o = n20122_o & n20123_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20125_o = n20121_o | n20124_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20126_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n20127_o = n20106_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n20128_o = n20126_o & n20127_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20129_o = n20125_o | n20128_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20130_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n20131_o = n20106_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n20132_o = n20130_o & n20131_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20133_o = n20129_o | n20132_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20134_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n20135_o = n20106_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n20136_o = n20134_o & n20135_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20137_o = n20133_o | n20136_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20138_o = ~n20137_o;
  /* vlm5030_gl.vhd:2281:16  */
  assign n20139_o = ~n20138_o;
  /* vlm5030_gl.vhd:2282:31  */
  assign n20141_o = aq[11];
  /* vlm5030_gl.vhd:2282:36  */
  assign n20142_o = {n20141_o, random};
  /* vlm5030_gl.vhd:2282:55  */
  assign n20144_o = {n20142_o, 1'b0};
  /* vlm5030_gl.vhd:2282:68  */
  assign n20146_o = {n20144_o, 1'b0};
  /* vlm5030_gl.vhd:2282:82  */
  assign n20147_o = {n20146_o, xromdo7nq};
  /* vlm5030_gl.vhd:2282:96  */
  assign n20149_o = {n20147_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n20155_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n20156_o = n20149_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n20157_o = n20155_o & n20156_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20159_o = 1'b0 | n20157_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20161_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n20162_o = n20149_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n20163_o = n20161_o & n20162_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20164_o = n20159_o | n20163_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20165_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n20166_o = n20149_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n20167_o = n20165_o & n20166_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20168_o = n20164_o | n20167_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20169_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n20170_o = n20149_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n20171_o = n20169_o & n20170_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20172_o = n20168_o | n20171_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20173_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n20174_o = n20149_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n20175_o = n20173_o & n20174_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20176_o = n20172_o | n20175_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20177_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n20178_o = n20149_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n20179_o = n20177_o & n20178_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20180_o = n20176_o | n20179_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20181_o = ~n20180_o;
  /* vlm5030_gl.vhd:2282:16  */
  assign n20182_o = ~n20181_o;
  /* vlm5030_gl.vhd:2283:31  */
  assign n20184_o = aq[12];
  /* vlm5030_gl.vhd:2283:49  */
  assign n20185_o = ieaddrreg[10];
  /* vlm5030_gl.vhd:2283:36  */
  assign n20186_o = {n20184_o, n20185_o};
  /* vlm5030_gl.vhd:2283:55  */
  assign n20188_o = {n20186_o, 1'b0};
  /* vlm5030_gl.vhd:2283:77  */
  assign n20189_o = nie[10];
  /* vlm5030_gl.vhd:2283:70  */
  assign n20190_o = ~n20189_o;
  /* vlm5030_gl.vhd:2283:68  */
  assign n20191_o = {n20188_o, n20190_o};
  /* vlm5030_gl.vhd:2283:91  */
  assign n20192_o = fsromdo[13];
  /* vlm5030_gl.vhd:2283:82  */
  assign n20193_o = {n20191_o, n20192_o};
  /* vlm5030_gl.vhd:2283:96  */
  assign n20195_o = {n20193_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n20201_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n20202_o = n20195_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n20203_o = n20201_o & n20202_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20205_o = 1'b0 | n20203_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20207_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n20208_o = n20195_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n20209_o = n20207_o & n20208_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20210_o = n20205_o | n20209_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20211_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n20212_o = n20195_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n20213_o = n20211_o & n20212_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20214_o = n20210_o | n20213_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20215_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n20216_o = n20195_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n20217_o = n20215_o & n20216_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20218_o = n20214_o | n20217_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20219_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n20220_o = n20195_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n20221_o = n20219_o & n20220_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20222_o = n20218_o | n20221_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20223_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n20224_o = n20195_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n20225_o = n20223_o & n20224_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20226_o = n20222_o | n20225_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20227_o = ~n20226_o;
  /* vlm5030_gl.vhd:2283:16  */
  assign n20228_o = ~n20227_o;
  /* vlm5030_gl.vhd:2284:31  */
  assign n20230_o = aq[13];
  /* vlm5030_gl.vhd:2284:49  */
  assign n20231_o = ieaddrreg[11];
  /* vlm5030_gl.vhd:2284:36  */
  assign n20232_o = {n20230_o, n20231_o};
  /* vlm5030_gl.vhd:2284:55  */
  assign n20234_o = {n20232_o, 1'b0};
  /* vlm5030_gl.vhd:2284:77  */
  assign n20235_o = nie[11];
  /* vlm5030_gl.vhd:2284:70  */
  assign n20236_o = ~n20235_o;
  /* vlm5030_gl.vhd:2284:68  */
  assign n20237_o = {n20234_o, n20236_o};
  /* vlm5030_gl.vhd:2284:82  */
  assign n20238_o = {n20237_o, vcufinal12};
  /* vlm5030_gl.vhd:2284:96  */
  assign n20240_o = {n20238_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n20246_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n20247_o = n20240_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n20248_o = n20246_o & n20247_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20250_o = 1'b0 | n20248_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20252_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n20253_o = n20240_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n20254_o = n20252_o & n20253_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20255_o = n20250_o | n20254_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20256_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n20257_o = n20240_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n20258_o = n20256_o & n20257_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20259_o = n20255_o | n20258_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20260_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n20261_o = n20240_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n20262_o = n20260_o & n20261_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20263_o = n20259_o | n20262_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20264_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n20265_o = n20240_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n20266_o = n20264_o & n20265_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20267_o = n20263_o | n20266_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20268_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n20269_o = n20240_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n20270_o = n20268_o & n20269_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20271_o = n20267_o | n20270_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20272_o = ~n20271_o;
  /* vlm5030_gl.vhd:2284:16  */
  assign n20273_o = ~n20272_o;
  /* vlm5030_gl.vhd:2285:31  */
  assign n20275_o = aq[14];
  /* vlm5030_gl.vhd:2285:36  */
  assign n20277_o = {n20275_o, 1'b0};
  /* vlm5030_gl.vhd:2285:55  */
  assign n20279_o = {n20277_o, 1'b0};
  /* vlm5030_gl.vhd:2285:68  */
  assign n20281_o = {n20279_o, 1'b0};
  /* vlm5030_gl.vhd:2285:82  */
  assign n20282_o = {n20281_o, cntdn0};
  /* vlm5030_gl.vhd:2285:96  */
  assign n20284_o = {n20282_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n20290_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n20291_o = n20284_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n20292_o = n20290_o & n20291_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20294_o = 1'b0 | n20292_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20296_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n20297_o = n20284_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n20298_o = n20296_o & n20297_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20299_o = n20294_o | n20298_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20300_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n20301_o = n20284_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n20302_o = n20300_o & n20301_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20303_o = n20299_o | n20302_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20304_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n20305_o = n20284_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n20306_o = n20304_o & n20305_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20307_o = n20303_o | n20306_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20308_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n20309_o = n20284_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n20310_o = n20308_o & n20309_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20311_o = n20307_o | n20310_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20312_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n20313_o = n20284_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n20314_o = n20312_o & n20313_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20315_o = n20311_o | n20314_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20316_o = ~n20315_o;
  /* vlm5030_gl.vhd:2285:16  */
  assign n20317_o = ~n20316_o;
  /* vlm5030_gl.vhd:2286:31  */
  assign n20319_o = aq[15];
  /* vlm5030_gl.vhd:2286:36  */
  assign n20321_o = {n20319_o, 1'b0};
  /* vlm5030_gl.vhd:2286:55  */
  assign n20323_o = {n20321_o, 1'b0};
  /* vlm5030_gl.vhd:2286:68  */
  assign n20325_o = {n20323_o, 1'b0};
  /* vlm5030_gl.vhd:2286:82  */
  assign n20327_o = {n20325_o, 1'b0};
  /* vlm5030_gl.vhd:2286:96  */
  assign n20329_o = {n20327_o, 1'b0};
  /* vlm5030_pack.vhd:50:26  */
  assign n20335_o = abus_block_wl[5];
  /* vlm5030_pack.vhd:50:39  */
  assign n20336_o = n20329_o[5];
  /* vlm5030_pack.vhd:50:32  */
  assign n20337_o = n20335_o & n20336_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20339_o = 1'b0 | n20337_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20341_o = abus_block_wl[4];
  /* vlm5030_pack.vhd:50:39  */
  assign n20342_o = n20329_o[4];
  /* vlm5030_pack.vhd:50:32  */
  assign n20343_o = n20341_o & n20342_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20344_o = n20339_o | n20343_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20345_o = abus_block_wl[3];
  /* vlm5030_pack.vhd:50:39  */
  assign n20346_o = n20329_o[3];
  /* vlm5030_pack.vhd:50:32  */
  assign n20347_o = n20345_o & n20346_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20348_o = n20344_o | n20347_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20349_o = abus_block_wl[2];
  /* vlm5030_pack.vhd:50:39  */
  assign n20350_o = n20329_o[2];
  /* vlm5030_pack.vhd:50:32  */
  assign n20351_o = n20349_o & n20350_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20352_o = n20348_o | n20351_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20353_o = abus_block_wl[1];
  /* vlm5030_pack.vhd:50:39  */
  assign n20354_o = n20329_o[1];
  /* vlm5030_pack.vhd:50:32  */
  assign n20355_o = n20353_o & n20354_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20356_o = n20352_o | n20355_o;
  /* vlm5030_pack.vhd:50:26  */
  assign n20357_o = abus_block_wl[0];
  /* vlm5030_pack.vhd:50:39  */
  assign n20358_o = n20329_o[0];
  /* vlm5030_pack.vhd:50:32  */
  assign n20359_o = n20357_o & n20358_o;
  /* vlm5030_pack.vhd:50:20  */
  assign n20360_o = n20356_o | n20359_o;
  /* vlm5030_pack.vhd:52:12  */
  assign n20361_o = ~n20360_o;
  /* vlm5030_gl.vhd:2286:16  */
  assign n20362_o = ~n20361_o;
  /* vlm5030_gl.vhd:2291:23  */
  assign n20363_o = ieaddrreg[9:0];
  /* vlm5030_gl.vhd:2291:53  */
  assign n20364_o = ~tstenie2dac;
  /* vlm5030_gl.vhd:2291:36  */
  assign n20365_o = n20364_o ? n20363_o : n20367_o;
  /* vlm5030_gl.vhd:2292:21  */
  assign n20366_o = nie[9:0];
  /* vlm5030_gl.vhd:2292:14  */
  assign n20367_o = ~n20366_o;
  /* vlm5030_gl.vhd:2294:12  */
  assign n20368_o = ~nbsy;
  /* vlm5030_gl.vhd:2296:13  */
  assign n20369_o = ~me;
  /* vlm5030_gl.vhd:2298:3  */
  vlm5030_delay_21 mte_delay_b (
    .i_clk_base(n20370_o),
    .i_clk_val(n20371_o),
    .i_clk_rise(n20372_o),
    .i_clk_fall(n20373_o),
    .i_in(n20374_o),
    .o_out(mte_delay_b_o_out));
  assign n20370_o = osc[0];
  assign n20371_o = osc[1];
  assign n20372_o = osc[2];
  assign n20373_o = osc[3];
  /* vlm5030_gl.vhd:2305:22  */
  assign n20374_o = xromdo[35];
  assign n20376_o = n8_o[1];
  assign n20377_o = clk2[1];
  /* vlm5030_gl.vhd:452:7  */
  assign n20378_o = n253_o ? n258_o : n20377_o;
  /* vlm5030_gl.vhd:452:7  */
  always @(posedge n251_o)
    n20379_q <= n20378_o;
  initial
    n20379_q = n20376_o;
  /* vlm5030_gl.vhd:452:7  */
  assign n20380_o = {n275_o, n263_o, n20379_q, n243_o};
  assign n20381_o = {n204_o, n203_o, n205_o};
  /* vlm5030_gl.vhd:495:7  */
  assign n20382_o = n305_o ? n308_o : clk2divq;
  /* vlm5030_gl.vhd:495:7  */
  always @(posedge n303_o)
    n20383_q <= n20382_o;
  initial
    n20383_q = 11'b00000000000;
  /* vlm5030_gl.vhd:662:9  */
  assign n20384_o = n2034_o ? n2058_o : xromdo7nq;
  /* vlm5030_gl.vhd:662:9  */
  always @(posedge n2032_o)
    n20385_q <= n20384_o;
  initial
    n20385_q = 1'b0;
  /* vlm5030_gl.vhd:854:7  */
  assign n20386_o = n5123_o ? n5127_o : dinalq;
  /* vlm5030_gl.vhd:854:7  */
  always @(posedge n5121_o or posedge clrdinal)
    if (clrdinal)
      n20387_q <= 8'b00000000;
    else
      n20387_q <= n20386_o;
  /* vlm5030_gl.vhd:875:7  */
  assign n20388_o = n5154_o ? n5165_o : aq;
  /* vlm5030_gl.vhd:875:7  */
  always @(posedge n5152_o)
    n20389_q <= n20388_o;
  /* vlm5030_gl.vhd:875:7  */
  assign n20390_o = {1'b0, n5861_o};
  assign n20391_o = {n15092_o, n15048_o, n15004_o, n14959_o, n14915_o, n14870_o, n14825_o, n14780_o, n14735_o, n14690_o};
  assign n20392_o = {n19489_o, n19447_o, n19405_o, n19363_o, n19318_o, n19273_o, n19228_o, n19183_o, n19138_o, n19093_o, n19048_o, n19003_o};
  /* vlm5030_gl.vhd:1609:7  */
  assign n20393_o = idlat_block_idlaten ? n15140_o : idlat;
  /* vlm5030_gl.vhd:1609:7  */
  always @(posedge n15138_o)
    n20394_q <= n20393_o;
  /* vlm5030_gl.vhd:1609:7  */
  assign n20395_o = {n18804_o, n18801_o, n18798_o, n18795_o, n18792_o, n18789_o, n18786_o, n18783_o, n18780_o, n18777_o, n18774_o, n18771_o};
  /* vlm5030_gl.vhd:2105:7  */
  assign n20396_o = n18901_o ? n18903_o : ieaddrreg;
  /* vlm5030_gl.vhd:2105:7  */
  always @(posedge n18899_o)
    n20397_q <= n20396_o;
  /* vlm5030_gl.vhd:2105:7  */
  assign n20398_o = {n20362_o, n20317_o, n20273_o, n20228_o, n20182_o, n20139_o, n20096_o, n20048_o, n20001_o, n19954_o, n19907_o, n19860_o, n19813_o, n19766_o, n19719_o, n19672_o};
  /* vlm5030_gl.vhd:1662:25  */
  reg [9:0] mem_block_mem0[9:0] ; // memory
  initial begin
    mem_block_mem0[9] = 10'b0000000000;
    mem_block_mem0[8] = 10'b0000000000;
    mem_block_mem0[7] = 10'b0000000000;
    mem_block_mem0[6] = 10'b0000000000;
    mem_block_mem0[5] = 10'b0000000000;
    mem_block_mem0[4] = 10'b0000000000;
    mem_block_mem0[3] = 10'b0000000000;
    mem_block_mem0[2] = 10'b0000000000;
    mem_block_mem0[1] = 10'b0000000000;
    mem_block_mem0[0] = 10'b0000000000;
    end
  assign n20400_data = mem_block_mem0[n15219_o];
  always @(posedge n15205_o)
    if (n15216_o)
      mem_block_mem0[n15210_o] <= nid;
  /* vlm5030_gl.vhd:1662:25  */
  /* vlm5030_gl.vhd:1655:18  */
  /* vlm5030_gl.vhd:1684:27  */
  reg [11:0] mem_block_mem1[9:0] ; // memory
  initial begin
    mem_block_mem1[9] = 12'b000000000000;
    mem_block_mem1[8] = 12'b000000000000;
    mem_block_mem1[7] = 12'b000000000000;
    mem_block_mem1[6] = 12'b000000000000;
    mem_block_mem1[5] = 12'b000000000000;
    mem_block_mem1[4] = 12'b000000000000;
    mem_block_mem1[3] = 12'b000000000000;
    mem_block_mem1[2] = 12'b000000000000;
    mem_block_mem1[1] = 12'b000000000000;
    mem_block_mem1[0] = 12'b000000000000;
    end
  assign n20403_data = mem_block_mem1[n15264_o];
  always @(posedge n15250_o)
    if (n15261_o)
      mem_block_mem1[n15255_o] <= nie;
  /* vlm5030_gl.vhd:1684:27  */
  /* vlm5030_gl.vhd:1677:18  */
  /* vlm5030_gl.vhd:1705:27  */
  reg [11:0] mem_block_mem2[8:0] ; // memory
  initial begin
    mem_block_mem2[8] = 12'b000000000000;
    mem_block_mem2[7] = 12'b000000000000;
    mem_block_mem2[6] = 12'b000000000000;
    mem_block_mem2[5] = 12'b000000000000;
    mem_block_mem2[4] = 12'b000000000000;
    mem_block_mem2[3] = 12'b000000000000;
    mem_block_mem2[2] = 12'b000000000000;
    mem_block_mem2[1] = 12'b000000000000;
    mem_block_mem2[0] = 12'b000000000000;
    end
  assign n20406_data = mem_block_mem2[n15309_o];
  always @(posedge n15295_o)
    if (n15306_o)
      mem_block_mem2[n15300_o] <= nie;
  /* vlm5030_gl.vhd:1705:27  */
  /* vlm5030_gl.vhd:1698:18  */
  /* vlm5030_gl.vhd:1219:9  */
  assign n20408_o = n5868_o[4];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20409_o = ~n20408_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20410_o = n5868_o[3];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20411_o = ~n20410_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20412_o = n20409_o & n20411_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20413_o = n20409_o & n20410_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20414_o = n20408_o & n20411_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20415_o = n20408_o & n20410_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20416_o = n5868_o[2];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20417_o = ~n20416_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20418_o = n20412_o & n20417_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20419_o = n20412_o & n20416_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20420_o = n20413_o & n20417_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20421_o = n20413_o & n20416_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20422_o = n20414_o & n20417_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20423_o = n20414_o & n20416_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20424_o = n20415_o & n20417_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20425_o = n20415_o & n20416_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20426_o = n5868_o[1];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20427_o = ~n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20428_o = n20418_o & n20427_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20429_o = n20418_o & n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20430_o = n20419_o & n20427_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20431_o = n20419_o & n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20432_o = n20420_o & n20427_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20433_o = n20420_o & n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20434_o = n20421_o & n20427_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20435_o = n20421_o & n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20436_o = n20422_o & n20427_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20437_o = n20422_o & n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20438_o = n20423_o & n20427_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20439_o = n20423_o & n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20440_o = n20424_o & n20427_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20441_o = n20424_o & n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20442_o = n20425_o & n20427_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20443_o = n20425_o & n20426_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20444_o = n5868_o[0];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20445_o = ~n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20446_o = n20428_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20447_o = n20428_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20448_o = n20429_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20449_o = n20429_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20450_o = n20430_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20451_o = n20430_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20452_o = n20431_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20453_o = n20431_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20454_o = n20432_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20455_o = n20432_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20456_o = n20433_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20457_o = n20433_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20458_o = n20434_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20459_o = n20434_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20460_o = n20435_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20461_o = n20435_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20462_o = n20436_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20463_o = n20436_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20464_o = n20437_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20465_o = n20437_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20466_o = n20438_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20467_o = n20438_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20468_o = n20439_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20469_o = n20439_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20470_o = n20440_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20471_o = n20440_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20472_o = n20441_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20473_o = n20441_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20474_o = n20442_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20475_o = n20442_o & n20444_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20476_o = n20443_o & n20445_o;
  /* vlm5030_gl.vhd:1219:9  */
  assign n20477_o = n20443_o & n20444_o;
  assign n20478_o = n5870_o[0];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20479_o = n20446_o ? 1'b1 : n20478_o;
  assign n20480_o = n5870_o[1];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20481_o = n20447_o ? 1'b1 : n20480_o;
  assign n20482_o = n5870_o[2];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20483_o = n20448_o ? 1'b1 : n20482_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20484_o = n5870_o[3];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20485_o = n20449_o ? 1'b1 : n20484_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20486_o = n5870_o[4];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20487_o = n20450_o ? 1'b1 : n20486_o;
  /* vlm5030_pack.vhd:46:14  */
  assign n20488_o = n5870_o[5];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20489_o = n20451_o ? 1'b1 : n20488_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20490_o = n5870_o[6];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20491_o = n20452_o ? 1'b1 : n20490_o;
  assign n20492_o = n5870_o[7];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20493_o = n20453_o ? 1'b1 : n20492_o;
  assign n20494_o = n5870_o[8];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20495_o = n20454_o ? 1'b1 : n20494_o;
  assign n20496_o = n5870_o[9];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20497_o = n20455_o ? 1'b1 : n20496_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20498_o = n5870_o[10];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20499_o = n20456_o ? 1'b1 : n20498_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20500_o = n5870_o[11];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20501_o = n20457_o ? 1'b1 : n20500_o;
  /* vlm5030_pack.vhd:46:14  */
  assign n20502_o = n5870_o[12];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20503_o = n20458_o ? 1'b1 : n20502_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20504_o = n5870_o[13];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20505_o = n20459_o ? 1'b1 : n20504_o;
  assign n20506_o = n5870_o[14];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20507_o = n20460_o ? 1'b1 : n20506_o;
  assign n20508_o = n5870_o[15];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20509_o = n20461_o ? 1'b1 : n20508_o;
  assign n20510_o = n5870_o[16];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20511_o = n20462_o ? 1'b1 : n20510_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20512_o = n5870_o[17];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20513_o = n20463_o ? 1'b1 : n20512_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20514_o = n5870_o[18];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20515_o = n20464_o ? 1'b1 : n20514_o;
  /* vlm5030_pack.vhd:46:14  */
  assign n20516_o = n5870_o[19];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20517_o = n20465_o ? 1'b1 : n20516_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20518_o = n5870_o[20];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20519_o = n20466_o ? 1'b1 : n20518_o;
  assign n20520_o = n5870_o[21];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20521_o = n20467_o ? 1'b1 : n20520_o;
  assign n20522_o = n5870_o[22];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20523_o = n20468_o ? 1'b1 : n20522_o;
  assign n20524_o = n5870_o[23];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20525_o = n20469_o ? 1'b1 : n20524_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20526_o = n5870_o[24];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20527_o = n20470_o ? 1'b1 : n20526_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20528_o = n5870_o[25];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20529_o = n20471_o ? 1'b1 : n20528_o;
  /* vlm5030_pack.vhd:46:14  */
  assign n20530_o = n5870_o[26];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20531_o = n20472_o ? 1'b1 : n20530_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20532_o = n5870_o[27];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20533_o = n20473_o ? 1'b1 : n20532_o;
  assign n20534_o = n5870_o[28];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20535_o = n20474_o ? 1'b1 : n20534_o;
  assign n20536_o = n5870_o[29];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20537_o = n20475_o ? 1'b1 : n20536_o;
  assign n20538_o = n5870_o[30];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20539_o = n20476_o ? 1'b1 : n20538_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20540_o = n5870_o[31];
  /* vlm5030_gl.vhd:1219:9  */
  assign n20541_o = n20477_o ? 1'b1 : n20540_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20542_o = {n20541_o, n20539_o, n20537_o, n20535_o, n20533_o, n20531_o, n20529_o, n20527_o, n20525_o, n20523_o, n20521_o, n20519_o, n20517_o, n20515_o, n20513_o, n20511_o, n20509_o, n20507_o, n20505_o, n20503_o, n20501_o, n20499_o, n20497_o, n20495_o, n20493_o, n20491_o, n20489_o, n20487_o, n20485_o, n20483_o, n20481_o, n20479_o};
  /* vlm5030_gl.vhd:1417:9  */
  assign n20543_o = n12790_o[3];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20544_o = ~n20543_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20545_o = n12790_o[2];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20546_o = ~n20545_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20547_o = n20544_o & n20546_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20548_o = n20544_o & n20545_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20549_o = n20543_o & n20546_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20550_o = n12790_o[1];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20551_o = ~n20550_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20552_o = n20547_o & n20551_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20553_o = n20547_o & n20550_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20554_o = n20548_o & n20551_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20555_o = n20548_o & n20550_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20556_o = n20549_o & n20551_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20557_o = n20549_o & n20550_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20558_o = n12790_o[0];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20559_o = ~n20558_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20560_o = n20552_o & n20559_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20561_o = n20552_o & n20558_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20562_o = n20553_o & n20559_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20563_o = n20553_o & n20558_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20564_o = n20554_o & n20559_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20565_o = n20554_o & n20558_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20566_o = n20555_o & n20559_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20567_o = n20555_o & n20558_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20568_o = n20556_o & n20559_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20569_o = n20556_o & n20558_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20570_o = n20557_o & n20559_o;
  /* vlm5030_gl.vhd:1417:9  */
  assign n20571_o = n20557_o & n20558_o;
  /* vlm5030_pack.vhd:26:13  */
  assign n20572_o = n12792_o[0];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20573_o = n20560_o ? 1'b1 : n20572_o;
  /* clock_functions_pack.vhd:65:34  */
  assign n20574_o = n12792_o[1];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20575_o = n20561_o ? 1'b1 : n20574_o;
  /* clock_functions_pack.vhd:35:12  */
  assign n20576_o = n12792_o[2];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20577_o = n20562_o ? 1'b1 : n20576_o;
  /* clock_functions_pack.vhd:35:12  */
  assign n20578_o = n12792_o[3];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20579_o = n20563_o ? 1'b1 : n20578_o;
  assign n20580_o = n12792_o[4];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20581_o = n20564_o ? 1'b1 : n20580_o;
  assign n20582_o = n12792_o[5];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20583_o = n20565_o ? 1'b1 : n20582_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20584_o = n12792_o[6];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20585_o = n20566_o ? 1'b1 : n20584_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20586_o = n12792_o[7];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20587_o = n20567_o ? 1'b1 : n20586_o;
  /* vlm5030_pack.vhd:46:14  */
  assign n20588_o = n12792_o[8];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20589_o = n20568_o ? 1'b1 : n20588_o;
  /* vlm5030_pack.vhd:27:13  */
  assign n20590_o = n12792_o[9];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20591_o = n20569_o ? 1'b1 : n20590_o;
  assign n20592_o = n12792_o[10];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20593_o = n20570_o ? 1'b1 : n20592_o;
  assign n20594_o = n12792_o[11];
  /* vlm5030_gl.vhd:1417:9  */
  assign n20595_o = n20571_o ? 1'b1 : n20594_o;
  assign n20596_o = {n20595_o, n20593_o, n20591_o, n20589_o, n20587_o, n20585_o, n20583_o, n20581_o, n20579_o, n20577_o, n20575_o, n20573_o};
endmodule

/* verilator lint_on UNOPTFLAT */