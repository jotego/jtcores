localparam [8:0]
    V_START  = 9'h100,
    VCNT_END = 9'h007,
    VB_START = 9'h000,
    VB_END   = 9'h120,
    VS_START = 9'h108,
    VS_END   = 9'h110;
