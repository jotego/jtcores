`timescale 1ns/1ps

module jtgng(
);



endmodule // jtgng