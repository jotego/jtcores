-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0b94",
     9 => x"ec080b0b",
    10 => x"0b94f008",
    11 => x"0b0b0b94",
    12 => x"f4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"94f40c0b",
    16 => x"0b0b94f0",
    17 => x"0c0b0b0b",
    18 => x"94ec0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0b94b8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"94ec7099",
    57 => x"c4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"81f70402",
    62 => x"e8050d83",
    63 => x"8b2d840b",
    64 => x"ec0c8ae5",
    65 => x"2d94ec08",
    66 => x"5394ec08",
    67 => x"802e80f2",
    68 => x"38850bec",
    69 => x"0c94c852",
    70 => x"94fc5191",
    71 => x"8d2d94ec",
    72 => x"08802e80",
    73 => x"d2389580",
    74 => x"08ff1154",
    75 => x"5572802e",
    76 => x"88387281",
    77 => x"2a5382ad",
    78 => x"04807525",
    79 => x"ba38958c",
    80 => x"5294fc51",
    81 => x"93c32d94",
    82 => x"ec08802e",
    83 => x"9a38958c",
    84 => x"5683fc54",
    85 => x"75708405",
    86 => x"5708e80c",
    87 => x"fc145473",
    88 => x"8025f138",
    89 => x"82ea0484",
    90 => x"805594fc",
    91 => x"5193962d",
    92 => x"fc801555",
    93 => x"82b90495",
    94 => x"8008f80c",
    95 => x"840bec0c",
    96 => x"80537294",
    97 => x"ec0c0298",
    98 => x"050d0481",
    99 => x"0bffb00c",
   100 => x"0402f405",
   101 => x"0dd45281",
   102 => x"ff720c71",
   103 => x"085381ff",
   104 => x"720c7288",
   105 => x"2b83fe80",
   106 => x"06720870",
   107 => x"81ff0651",
   108 => x"525381ff",
   109 => x"720c7271",
   110 => x"07882b72",
   111 => x"087081ff",
   112 => x"06515253",
   113 => x"81ff720c",
   114 => x"72710788",
   115 => x"2b720870",
   116 => x"81ff0672",
   117 => x"0794ec0c",
   118 => x"5253028c",
   119 => x"050d0402",
   120 => x"f4050d74",
   121 => x"767181ff",
   122 => x"06d40c53",
   123 => x"53958808",
   124 => x"85387189",
   125 => x"2b527198",
   126 => x"2ad40c71",
   127 => x"902a7081",
   128 => x"ff06d40c",
   129 => x"5171882a",
   130 => x"7081ff06",
   131 => x"d40c5171",
   132 => x"81ff06d4",
   133 => x"0c72902a",
   134 => x"7081ff06",
   135 => x"d40c51d4",
   136 => x"087081ff",
   137 => x"06515182",
   138 => x"b8bf5270",
   139 => x"81ff2e09",
   140 => x"81069438",
   141 => x"81ff0bd4",
   142 => x"0cd40870",
   143 => x"81ff06ff",
   144 => x"14545151",
   145 => x"71e53870",
   146 => x"94ec0c02",
   147 => x"8c050d04",
   148 => x"02fc050d",
   149 => x"81c75181",
   150 => x"ff0bd40c",
   151 => x"ff115170",
   152 => x"8025f438",
   153 => x"0284050d",
   154 => x"0402f405",
   155 => x"0d81ff0b",
   156 => x"d40c9353",
   157 => x"805287fc",
   158 => x"80c15183",
   159 => x"df2d94ec",
   160 => x"088b3881",
   161 => x"ff0bd40c",
   162 => x"81538596",
   163 => x"0484d02d",
   164 => x"ff135372",
   165 => x"df387294",
   166 => x"ec0c028c",
   167 => x"050d0402",
   168 => x"ec050d81",
   169 => x"0b95880c",
   170 => x"8454d008",
   171 => x"708f2a70",
   172 => x"81065151",
   173 => x"5372f338",
   174 => x"72d00c84",
   175 => x"d02dd008",
   176 => x"708f2a70",
   177 => x"81065151",
   178 => x"5372f338",
   179 => x"810bd00c",
   180 => x"b1538052",
   181 => x"84d480c0",
   182 => x"5183df2d",
   183 => x"94ec0881",
   184 => x"2e933872",
   185 => x"822ebd38",
   186 => x"ff135372",
   187 => x"e538ff14",
   188 => x"5473ffb6",
   189 => x"3884d02d",
   190 => x"83aa5284",
   191 => x"9c80c851",
   192 => x"83df2d94",
   193 => x"ec08812e",
   194 => x"09810692",
   195 => x"3883912d",
   196 => x"94ec0883",
   197 => x"ffff0653",
   198 => x"7283aa2e",
   199 => x"913884e9",
   200 => x"2d86a904",
   201 => x"805387f7",
   202 => x"04805487",
   203 => x"c90481ff",
   204 => x"0bd40cb1",
   205 => x"5484d02d",
   206 => x"8fcf5380",
   207 => x"5287fc80",
   208 => x"f75183df",
   209 => x"2d94ec08",
   210 => x"5594ec08",
   211 => x"812e0981",
   212 => x"069b3881",
   213 => x"ff0bd40c",
   214 => x"820a5284",
   215 => x"9c80e951",
   216 => x"83df2d94",
   217 => x"ec08802e",
   218 => x"8d3884d0",
   219 => x"2dff1353",
   220 => x"72c93887",
   221 => x"bc0481ff",
   222 => x"0bd40c94",
   223 => x"ec085287",
   224 => x"fc80fa51",
   225 => x"83df2d94",
   226 => x"ec08b138",
   227 => x"81ff0bd4",
   228 => x"0cd40853",
   229 => x"81ff0bd4",
   230 => x"0c81ff0b",
   231 => x"d40c81ff",
   232 => x"0bd40c81",
   233 => x"ff0bd40c",
   234 => x"72862a70",
   235 => x"81067656",
   236 => x"51537295",
   237 => x"3894ec08",
   238 => x"5487c904",
   239 => x"73822efe",
   240 => x"e838ff14",
   241 => x"5473feed",
   242 => x"38739588",
   243 => x"0c738b38",
   244 => x"815287fc",
   245 => x"80d05183",
   246 => x"df2d81ff",
   247 => x"0bd40cd0",
   248 => x"08708f2a",
   249 => x"70810651",
   250 => x"515372f3",
   251 => x"3872d00c",
   252 => x"81ff0bd4",
   253 => x"0c815372",
   254 => x"94ec0c02",
   255 => x"94050d04",
   256 => x"02e8050d",
   257 => x"78558056",
   258 => x"81ff0bd4",
   259 => x"0cd00870",
   260 => x"8f2a7081",
   261 => x"06515153",
   262 => x"72f33882",
   263 => x"810bd00c",
   264 => x"81ff0bd4",
   265 => x"0c775287",
   266 => x"fc80d151",
   267 => x"83df2d94",
   268 => x"ec0880d9",
   269 => x"3880dbc6",
   270 => x"df5481ff",
   271 => x"0bd40cd4",
   272 => x"087081ff",
   273 => x"06515372",
   274 => x"81fe2e09",
   275 => x"81069d38",
   276 => x"80ff5383",
   277 => x"912d94ec",
   278 => x"08757084",
   279 => x"05570cff",
   280 => x"13537280",
   281 => x"25ed3881",
   282 => x"5688f204",
   283 => x"ff145473",
   284 => x"c93881ff",
   285 => x"0bd40c81",
   286 => x"ff0bd40c",
   287 => x"d008708f",
   288 => x"2a708106",
   289 => x"51515372",
   290 => x"f33872d0",
   291 => x"0c7594ec",
   292 => x"0c029805",
   293 => x"0d0402e8",
   294 => x"050d7779",
   295 => x"7b585555",
   296 => x"80537276",
   297 => x"25a33874",
   298 => x"70810556",
   299 => x"80f52d74",
   300 => x"70810556",
   301 => x"80f52d52",
   302 => x"5271712e",
   303 => x"86388151",
   304 => x"89cb0481",
   305 => x"135389a2",
   306 => x"04805170",
   307 => x"94ec0c02",
   308 => x"98050d04",
   309 => x"02ec050d",
   310 => x"76557480",
   311 => x"2ebb389a",
   312 => x"1580e02d",
   313 => x"5194992d",
   314 => x"94ec0894",
   315 => x"ec0899b8",
   316 => x"0c94ec08",
   317 => x"54549994",
   318 => x"08802e99",
   319 => x"38941580",
   320 => x"e02d5194",
   321 => x"992d94ec",
   322 => x"08902b83",
   323 => x"fff00a06",
   324 => x"70750751",
   325 => x"537299b8",
   326 => x"0c99b808",
   327 => x"5372802e",
   328 => x"9938998c",
   329 => x"08fe1471",
   330 => x"2999a008",
   331 => x"0599bc0c",
   332 => x"70842b99",
   333 => x"980c548a",
   334 => x"e00499a4",
   335 => x"0899b80c",
   336 => x"99a80899",
   337 => x"bc0c9994",
   338 => x"08802e8a",
   339 => x"38998c08",
   340 => x"842b538a",
   341 => x"dc0499ac",
   342 => x"08842b53",
   343 => x"7299980c",
   344 => x"0294050d",
   345 => x"0402d805",
   346 => x"0d800b99",
   347 => x"940c8454",
   348 => x"859f2d94",
   349 => x"ec08802e",
   350 => x"9538958c",
   351 => x"52805188",
   352 => x"802d94ec",
   353 => x"08802e86",
   354 => x"38fe548b",
   355 => x"9604ff14",
   356 => x"54738024",
   357 => x"db387355",
   358 => x"73802e84",
   359 => x"f9388056",
   360 => x"810b99c0",
   361 => x"0c885394",
   362 => x"d45295c2",
   363 => x"5189962d",
   364 => x"94ec0876",
   365 => x"2e098106",
   366 => x"873894ec",
   367 => x"0899c00c",
   368 => x"885394e0",
   369 => x"5295de51",
   370 => x"89962d94",
   371 => x"ec088738",
   372 => x"94ec0899",
   373 => x"c00c99c0",
   374 => x"08802e80",
   375 => x"f63898d2",
   376 => x"0b80f52d",
   377 => x"98d30b80",
   378 => x"f52d7198",
   379 => x"2b71902b",
   380 => x"0798d40b",
   381 => x"80f52d70",
   382 => x"882b7207",
   383 => x"98d50b80",
   384 => x"f52d7107",
   385 => x"998a0b80",
   386 => x"f52d998b",
   387 => x"0b80f52d",
   388 => x"71882b07",
   389 => x"535f5452",
   390 => x"5a565755",
   391 => x"7381abaa",
   392 => x"2e098106",
   393 => x"8d387551",
   394 => x"93e92d94",
   395 => x"ec08568c",
   396 => x"bf048055",
   397 => x"7382d4d5",
   398 => x"2e098106",
   399 => x"83d83895",
   400 => x"8c527551",
   401 => x"88802d94",
   402 => x"ec085594",
   403 => x"ec08802e",
   404 => x"83c43888",
   405 => x"5394e052",
   406 => x"95de5189",
   407 => x"962d94ec",
   408 => x"08893881",
   409 => x"0b99940c",
   410 => x"8d830488",
   411 => x"5394d452",
   412 => x"95c25189",
   413 => x"962d8055",
   414 => x"94ec0875",
   415 => x"2e098106",
   416 => x"83943899",
   417 => x"8a0b80f5",
   418 => x"2d547380",
   419 => x"d52e0981",
   420 => x"0680ca38",
   421 => x"998b0b80",
   422 => x"f52d5473",
   423 => x"81aa2e09",
   424 => x"8106ba38",
   425 => x"800b958c",
   426 => x"0b80f52d",
   427 => x"56547481",
   428 => x"e92e8338",
   429 => x"81547481",
   430 => x"eb2e8c38",
   431 => x"80557375",
   432 => x"2e098106",
   433 => x"82d03895",
   434 => x"970b80f5",
   435 => x"2d55748d",
   436 => x"3895980b",
   437 => x"80f52d54",
   438 => x"73822e86",
   439 => x"38805590",
   440 => x"96049599",
   441 => x"0b80f52d",
   442 => x"70998c0c",
   443 => x"ff059990",
   444 => x"0c959a0b",
   445 => x"80f52d95",
   446 => x"9b0b80f5",
   447 => x"2d587605",
   448 => x"77828029",
   449 => x"0570999c",
   450 => x"0c959c0b",
   451 => x"80f52d70",
   452 => x"99b00c99",
   453 => x"94085957",
   454 => x"5876802e",
   455 => x"81a33888",
   456 => x"5394e052",
   457 => x"95de5189",
   458 => x"962d94ec",
   459 => x"0881e738",
   460 => x"998c0870",
   461 => x"842b9998",
   462 => x"0c7099ac",
   463 => x"0c95b10b",
   464 => x"80f52d95",
   465 => x"b00b80f5",
   466 => x"2d718280",
   467 => x"290595b2",
   468 => x"0b80f52d",
   469 => x"70848080",
   470 => x"291295b3",
   471 => x"0b80f52d",
   472 => x"7081800a",
   473 => x"29127099",
   474 => x"b40c99b0",
   475 => x"08712999",
   476 => x"9c080570",
   477 => x"99a00c95",
   478 => x"b90b80f5",
   479 => x"2d95b80b",
   480 => x"80f52d71",
   481 => x"82802905",
   482 => x"95ba0b80",
   483 => x"f52d7084",
   484 => x"80802912",
   485 => x"95bb0b80",
   486 => x"f52d7098",
   487 => x"2b81f00a",
   488 => x"06720570",
   489 => x"99a40cfe",
   490 => x"117e2977",
   491 => x"0599a80c",
   492 => x"52595243",
   493 => x"545e5152",
   494 => x"59525d57",
   495 => x"5957908f",
   496 => x"04959e0b",
   497 => x"80f52d95",
   498 => x"9d0b80f5",
   499 => x"2d718280",
   500 => x"29057099",
   501 => x"980c70a0",
   502 => x"2983ff05",
   503 => x"70892a70",
   504 => x"99ac0c95",
   505 => x"a30b80f5",
   506 => x"2d95a20b",
   507 => x"80f52d71",
   508 => x"82802905",
   509 => x"7099b40c",
   510 => x"7b71291e",
   511 => x"7099a80c",
   512 => x"7d99a40c",
   513 => x"730599a0",
   514 => x"0c555e51",
   515 => x"51555580",
   516 => x"5189d42d",
   517 => x"81557494",
   518 => x"ec0c02a8",
   519 => x"050d0402",
   520 => x"ec050d76",
   521 => x"70872c71",
   522 => x"80ff0655",
   523 => x"56549994",
   524 => x"088a3873",
   525 => x"882c7481",
   526 => x"ff065455",
   527 => x"958c5299",
   528 => x"9c081551",
   529 => x"88802d94",
   530 => x"ec085494",
   531 => x"ec08802e",
   532 => x"b3389994",
   533 => x"08802e98",
   534 => x"38728429",
   535 => x"958c0570",
   536 => x"08525393",
   537 => x"e92d94ec",
   538 => x"08f00a06",
   539 => x"53918204",
   540 => x"7210958c",
   541 => x"057080e0",
   542 => x"2d525394",
   543 => x"992d94ec",
   544 => x"08537254",
   545 => x"7394ec0c",
   546 => x"0294050d",
   547 => x"0402cc05",
   548 => x"0d7e605e",
   549 => x"5a800b99",
   550 => x"b80899bc",
   551 => x"08595c56",
   552 => x"80589998",
   553 => x"08782e81",
   554 => x"ae38778f",
   555 => x"06a01757",
   556 => x"54738f38",
   557 => x"958c5276",
   558 => x"51811757",
   559 => x"88802d95",
   560 => x"8c568076",
   561 => x"80f52d56",
   562 => x"5474742e",
   563 => x"83388154",
   564 => x"7481e52e",
   565 => x"80f63881",
   566 => x"70750655",
   567 => x"5c73802e",
   568 => x"80ea388b",
   569 => x"1680f52d",
   570 => x"98065978",
   571 => x"80de388b",
   572 => x"537c5275",
   573 => x"5189962d",
   574 => x"94ec0880",
   575 => x"cf389c16",
   576 => x"085193e9",
   577 => x"2d94ec08",
   578 => x"841b0c9a",
   579 => x"1680e02d",
   580 => x"5194992d",
   581 => x"94ec0894",
   582 => x"ec08881c",
   583 => x"0c94ec08",
   584 => x"55559994",
   585 => x"08802e98",
   586 => x"38941680",
   587 => x"e02d5194",
   588 => x"992d94ec",
   589 => x"08902b83",
   590 => x"fff00a06",
   591 => x"70165154",
   592 => x"73881b0c",
   593 => x"787a0c7b",
   594 => x"54938d04",
   595 => x"81185899",
   596 => x"98087826",
   597 => x"fed43899",
   598 => x"9408802e",
   599 => x"ae387a51",
   600 => x"909f2d94",
   601 => x"ec0894ec",
   602 => x"0880ffff",
   603 => x"fff80655",
   604 => x"5b7380ff",
   605 => x"fffff82e",
   606 => x"923894ec",
   607 => x"08fe0599",
   608 => x"8c082999",
   609 => x"a0080557",
   610 => x"91a00480",
   611 => x"547394ec",
   612 => x"0c02b405",
   613 => x"0d0402f4",
   614 => x"050d7470",
   615 => x"08810571",
   616 => x"0c700899",
   617 => x"90080653",
   618 => x"53718e38",
   619 => x"88130851",
   620 => x"909f2d94",
   621 => x"ec088814",
   622 => x"0c810b94",
   623 => x"ec0c028c",
   624 => x"050d0402",
   625 => x"f0050d75",
   626 => x"881108fe",
   627 => x"05998c08",
   628 => x"2999a008",
   629 => x"11720899",
   630 => x"90080605",
   631 => x"79555354",
   632 => x"5488802d",
   633 => x"0290050d",
   634 => x"0402f405",
   635 => x"0d747088",
   636 => x"2a83fe80",
   637 => x"06707298",
   638 => x"2a077288",
   639 => x"2b87fc80",
   640 => x"80067398",
   641 => x"2b81f00a",
   642 => x"06717307",
   643 => x"0794ec0c",
   644 => x"56515351",
   645 => x"028c050d",
   646 => x"0402f805",
   647 => x"0d028e05",
   648 => x"80f52d74",
   649 => x"882b0770",
   650 => x"83ffff06",
   651 => x"94ec0c51",
   652 => x"0288050d",
   653 => x"04000000",
   654 => x"00ffffff",
   655 => x"ff00ffff",
   656 => x"ffff00ff",
   657 => x"ffffff00",
   658 => x"4a54474e",
   659 => x"47202020",
   660 => x"524f4d00",
   661 => x"46415431",
   662 => x"36202020",
   663 => x"00000000",
   664 => x"46415433",
   665 => x"32202020",
   666 => x"00202020",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

