/*  This file is part of JT_GNG.
    JT_GNG program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT_GNG program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT_GNG.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 5-4-2021 */

module jtrumble_banks(
    input      [7:0] msb_addr,
    input      [7:0] lsb_addr,
    output reg [3:0] msb,
    output reg [3:0] lsb
);

always@(msb_addr)
    case( msb_addr )
          0: msb=4'h0;
          1: msb=4'h0;
          2: msb=4'h0;
          3: msb=4'h0;
          4: msb=4'h1;
          5: msb=4'h0;
          6: msb=4'h0;
          7: msb=4'h7;
          8: msb=4'h7;
          9: msb=4'h7;
         10: msb=4'h7;
         11: msb=4'h4;
         12: msb=4'h4;
         13: msb=4'h4;
         14: msb=4'h4;
         15: msb=4'h4;
         16: msb=4'h0;
         17: msb=4'h0;
         18: msb=4'h0;
         19: msb=4'h0;
         20: msb=4'h1;
         21: msb=4'h0;
         22: msb=4'h0;
         23: msb=4'h0;
         24: msb=4'h0;
         25: msb=4'h4;
         26: msb=4'h5;
         27: msb=4'h4;
         28: msb=4'h4;
         29: msb=4'h4;
         30: msb=4'h4;
         31: msb=4'h4;
         32: msb=4'h0;
         33: msb=4'h0;
         34: msb=4'h0;
         35: msb=4'h0;
         36: msb=4'h1;
         37: msb=4'h4;
         38: msb=4'h4;
         39: msb=4'h4;
         40: msb=4'h4;
         41: msb=4'h4;
         42: msb=4'h4;
         43: msb=4'h4;
         44: msb=4'h4;
         45: msb=4'h5;
         46: msb=4'h4;
         47: msb=4'h4;
         48: msb=4'h0;
         49: msb=4'h0;
         50: msb=4'h0;
         51: msb=4'h0;
         52: msb=4'h1;
         53: msb=4'h4;
         54: msb=4'h4;
         55: msb=4'h7;
         56: msb=4'h7;
         57: msb=4'h7;
         58: msb=4'h7;
         59: msb=4'h4;
         60: msb=4'h4;
         61: msb=4'h4;
         62: msb=4'h4;
         63: msb=4'h4;
         64: msb=4'h0;
         65: msb=4'h0;
         66: msb=4'h0;
         67: msb=4'h0;
         68: msb=4'h1;
         69: msb=4'h4;
         70: msb=4'h4;
         71: msb=4'h4;
         72: msb=4'h4;
         73: msb=4'h5;
         74: msb=4'h5;
         75: msb=4'h5;
         76: msb=4'h5;
         77: msb=4'h5;
         78: msb=4'h4;
         79: msb=4'h4;
         80: msb=4'h0;
         81: msb=4'h0;
         82: msb=4'h0;
         83: msb=4'h0;
         84: msb=4'h1;
         85: msb=4'h5;
         86: msb=4'h5;
         87: msb=4'h5;
         88: msb=4'h5;
         89: msb=4'h5;
         90: msb=4'h5;
         91: msb=4'h5;
         92: msb=4'h5;
         93: msb=4'h5;
         94: msb=4'h4;
         95: msb=4'h4;
         96: msb=4'h0;
         97: msb=4'h0;
         98: msb=4'h0;
         99: msb=4'h0;
        100: msb=4'h1;
        101: msb=4'h4;
        102: msb=4'h4;
        103: msb=4'h4;
        104: msb=4'h4;
        105: msb=4'h6;
        106: msb=4'h6;
        107: msb=4'h6;
        108: msb=4'h6;
        109: msb=4'h5;
        110: msb=4'h4;
        111: msb=4'h4;
        112: msb=4'h0;
        113: msb=4'h0;
        114: msb=4'h0;
        115: msb=4'h0;
        116: msb=4'h1;
        117: msb=4'h4;
        118: msb=4'h4;
        119: msb=4'h4;
        120: msb=4'h4;
        121: msb=4'h6;
        122: msb=4'h6;
        123: msb=4'h6;
        124: msb=4'h6;
        125: msb=4'h6;
        126: msb=4'h4;
        127: msb=4'h4;
        128: msb=4'h0;
        129: msb=4'h0;
        130: msb=4'h0;
        131: msb=4'h0;
        132: msb=4'h1;
        133: msb=4'h0;
        134: msb=4'h0;
        135: msb=4'h7;
        136: msb=4'h7;
        137: msb=4'h7;
        138: msb=4'h7;
        139: msb=4'h4;
        140: msb=4'h4;
        141: msb=4'h4;
        142: msb=4'h4;
        143: msb=4'h4;
        144: msb=4'h0;
        145: msb=4'h0;
        146: msb=4'h0;
        147: msb=4'h0;
        148: msb=4'h1;
        149: msb=4'h0;
        150: msb=4'h0;
        151: msb=4'h7;
        152: msb=4'h7;
        153: msb=4'h7;
        154: msb=4'h7;
        155: msb=4'h4;
        156: msb=4'h4;
        157: msb=4'h4;
        158: msb=4'h4;
        159: msb=4'h4;
        160: msb=4'h0;
        161: msb=4'h0;
        162: msb=4'h0;
        163: msb=4'h0;
        164: msb=4'h1;
        165: msb=4'h0;
        166: msb=4'h0;
        167: msb=4'h7;
        168: msb=4'h7;
        169: msb=4'h7;
        170: msb=4'h7;
        171: msb=4'h4;
        172: msb=4'h4;
        173: msb=4'h4;
        174: msb=4'h4;
        175: msb=4'h4;
        176: msb=4'h0;
        177: msb=4'h0;
        178: msb=4'h0;
        179: msb=4'h0;
        180: msb=4'h1;
        181: msb=4'h0;
        182: msb=4'h0;
        183: msb=4'h7;
        184: msb=4'h7;
        185: msb=4'h7;
        186: msb=4'h7;
        187: msb=4'h4;
        188: msb=4'h4;
        189: msb=4'h4;
        190: msb=4'h4;
        191: msb=4'h4;
        192: msb=4'h0;
        193: msb=4'h0;
        194: msb=4'h0;
        195: msb=4'h0;
        196: msb=4'h1;
        197: msb=4'h0;
        198: msb=4'h0;
        199: msb=4'h7;
        200: msb=4'h7;
        201: msb=4'h7;
        202: msb=4'h7;
        203: msb=4'h4;
        204: msb=4'h4;
        205: msb=4'h4;
        206: msb=4'h4;
        207: msb=4'h4;
        208: msb=4'h0;
        209: msb=4'h0;
        210: msb=4'h0;
        211: msb=4'h0;
        212: msb=4'h1;
        213: msb=4'h0;
        214: msb=4'h0;
        215: msb=4'h7;
        216: msb=4'h7;
        217: msb=4'h7;
        218: msb=4'h7;
        219: msb=4'h4;
        220: msb=4'h4;
        221: msb=4'h4;
        222: msb=4'h4;
        223: msb=4'h4;
        224: msb=4'h0;
        225: msb=4'h0;
        226: msb=4'h0;
        227: msb=4'h0;
        228: msb=4'h1;
        229: msb=4'h0;
        230: msb=4'h0;
        231: msb=4'h7;
        232: msb=4'h7;
        233: msb=4'h7;
        234: msb=4'h7;
        235: msb=4'h4;
        236: msb=4'h4;
        237: msb=4'h4;
        238: msb=4'h4;
        239: msb=4'h4;
        240: msb=4'h0;
        241: msb=4'h0;
        242: msb=4'h0;
        243: msb=4'h0;
        244: msb=4'h1;
        245: msb=4'h0;
        246: msb=4'h0;
        247: msb=4'h7;
        248: msb=4'h7;
        249: msb=4'h7;
        250: msb=4'h7;
        251: msb=4'h4;
        252: msb=4'h4;
        253: msb=4'h4;
        254: msb=4'h4;
        255: msb=4'h4;
    endcase

always @(lsb_addr)
    case( lsb_addr )
          0: lsb=4'h0;
          1: lsb=4'h1;
          2: lsb=4'h4;
          3: lsb=4'h5;
          4: lsb=4'h0;
          5: lsb=4'h8;
          6: lsb=4'h9;
          7: lsb=4'hC;
          8: lsb=4'hD;
          9: lsb=4'hE;
         10: lsb=4'hF;
         11: lsb=4'hB;
         12: lsb=4'hE;
         13: lsb=4'hF;
         14: lsb=4'hC;
         15: lsb=4'hD;
         16: lsb=4'h0;
         17: lsb=4'h1;
         18: lsb=4'h4;
         19: lsb=4'h5;
         20: lsb=4'h0;
         21: lsb=4'h8;
         22: lsb=4'h9;
         23: lsb=4'h0;
         24: lsb=4'h1;
         25: lsb=4'h2;
         26: lsb=4'h3;
         27: lsb=4'hB;
         28: lsb=4'hE;
         29: lsb=4'hF;
         30: lsb=4'hC;
         31: lsb=4'hD;
         32: lsb=4'h0;
         33: lsb=4'h1;
         34: lsb=4'h4;
         35: lsb=4'h5;
         36: lsb=4'h0;
         37: lsb=4'h8;
         38: lsb=4'h9;
         39: lsb=4'h4;
         40: lsb=4'h5;
         41: lsb=4'h6;
         42: lsb=4'h7;
         43: lsb=4'hB;
         44: lsb=4'hE;
         45: lsb=4'hF;
         46: lsb=4'hC;
         47: lsb=4'hD;
         48: lsb=4'h0;
         49: lsb=4'h1;
         50: lsb=4'h4;
         51: lsb=4'h5;
         52: lsb=4'h0;
         53: lsb=4'h8;
         54: lsb=4'h9;
         55: lsb=4'h8;
         56: lsb=4'h9;
         57: lsb=4'hA;
         58: lsb=4'hB;
         59: lsb=4'hB;
         60: lsb=4'hE;
         61: lsb=4'hF;
         62: lsb=4'hC;
         63: lsb=4'hD;
         64: lsb=4'h0;
         65: lsb=4'h1;
         66: lsb=4'h4;
         67: lsb=4'h5;
         68: lsb=4'h0;
         69: lsb=4'h8;
         70: lsb=4'h9;
         71: lsb=4'hC;
         72: lsb=4'hD;
         73: lsb=4'hA;
         74: lsb=4'h6;
         75: lsb=4'hB;
         76: lsb=4'hE;
         77: lsb=4'hF;
         78: lsb=4'hC;
         79: lsb=4'hD;
         80: lsb=4'h0;
         81: lsb=4'h1;
         82: lsb=4'h4;
         83: lsb=4'h5;
         84: lsb=4'h0;
         85: lsb=4'h0;
         86: lsb=4'h1;
         87: lsb=4'h2;
         88: lsb=4'h3;
         89: lsb=4'h4;
         90: lsb=4'h5;
         91: lsb=4'h6;
         92: lsb=4'h7;
         93: lsb=4'h7;
         94: lsb=4'hC;
         95: lsb=4'hD;
         96: lsb=4'h0;
         97: lsb=4'h1;
         98: lsb=4'h4;
         99: lsb=4'h5;
        100: lsb=4'h0;
        101: lsb=4'h0;
        102: lsb=4'h1;
        103: lsb=4'h2;
        104: lsb=4'h3;
        105: lsb=4'h0;
        106: lsb=4'h1;
        107: lsb=4'h2;
        108: lsb=4'h3;
        109: lsb=4'h4;
        110: lsb=4'hC;
        111: lsb=4'hD;
        112: lsb=4'h0;
        113: lsb=4'h1;
        114: lsb=4'h4;
        115: lsb=4'h5;
        116: lsb=4'h0;
        117: lsb=4'h0;
        118: lsb=4'h1;
        119: lsb=4'h2;
        120: lsb=4'h3;
        121: lsb=4'h2;
        122: lsb=4'h3;
        123: lsb=4'h4;
        124: lsb=4'h5;
        125: lsb=4'h6;
        126: lsb=4'hC;
        127: lsb=4'hD;
        128: lsb=4'h0;
        129: lsb=4'h1;
        130: lsb=4'h4;
        131: lsb=4'h5;
        132: lsb=4'h0;
        133: lsb=4'h8;
        134: lsb=4'h9;
        135: lsb=4'hA;
        136: lsb=4'hB;
        137: lsb=4'hC;
        138: lsb=4'hD;
        139: lsb=4'hE;
        140: lsb=4'hF;
        141: lsb=4'h0;
        142: lsb=4'hC;
        143: lsb=4'hD;
        144: lsb=4'h0;
        145: lsb=4'h1;
        146: lsb=4'h4;
        147: lsb=4'h5;
        148: lsb=4'h0;
        149: lsb=4'h0;
        150: lsb=4'h1;
        151: lsb=4'h2;
        152: lsb=4'h3;
        153: lsb=4'h0;
        154: lsb=4'h1;
        155: lsb=4'h2;
        156: lsb=4'h3;
        157: lsb=4'h7;
        158: lsb=4'hC;
        159: lsb=4'hD;
        160: lsb=4'h0;
        161: lsb=4'h1;
        162: lsb=4'h4;
        163: lsb=4'h5;
        164: lsb=4'h0;
        165: lsb=4'h0;
        166: lsb=4'h1;
        167: lsb=4'h2;
        168: lsb=4'h3;
        169: lsb=4'h4;
        170: lsb=4'h5;
        171: lsb=4'h6;
        172: lsb=4'h7;
        173: lsb=4'h6;
        174: lsb=4'hC;
        175: lsb=4'hD;
        176: lsb=4'h0;
        177: lsb=4'h1;
        178: lsb=4'h4;
        179: lsb=4'h5;
        180: lsb=4'h0;
        181: lsb=4'h0;
        182: lsb=4'h1;
        183: lsb=4'h2;
        184: lsb=4'h3;
        185: lsb=4'h8;
        186: lsb=4'h9;
        187: lsb=4'hA;
        188: lsb=4'hB;
        189: lsb=4'h6;
        190: lsb=4'hC;
        191: lsb=4'hD;
        192: lsb=4'h0;
        193: lsb=4'h1;
        194: lsb=4'h4;
        195: lsb=4'h5;
        196: lsb=4'h0;
        197: lsb=4'h0;
        198: lsb=4'h1;
        199: lsb=4'h2;
        200: lsb=4'h3;
        201: lsb=4'hC;
        202: lsb=4'hD;
        203: lsb=4'hE;
        204: lsb=4'hF;
        205: lsb=4'h7;
        206: lsb=4'hC;
        207: lsb=4'hD;
        208: lsb=4'h0;
        209: lsb=4'h1;
        210: lsb=4'h4;
        211: lsb=4'h5;
        212: lsb=4'h0;
        213: lsb=4'h0;
        214: lsb=4'h1;
        215: lsb=4'h2;
        216: lsb=4'h3;
        217: lsb=4'h6;
        218: lsb=4'h7;
        219: lsb=4'h0;
        220: lsb=4'h1;
        221: lsb=4'h2;
        222: lsb=4'hC;
        223: lsb=4'hD;
        224: lsb=4'h0;
        225: lsb=4'h1;
        226: lsb=4'h4;
        227: lsb=4'h5;
        228: lsb=4'h0;
        229: lsb=4'h0;
        230: lsb=4'h1;
        231: lsb=4'h2;
        232: lsb=4'h3;
        233: lsb=4'h6;
        234: lsb=4'h7;
        235: lsb=4'h0;
        236: lsb=4'h1;
        237: lsb=4'h7;
        238: lsb=4'hC;
        239: lsb=4'hD;
        240: lsb=4'h0;
        241: lsb=4'h1;
        242: lsb=4'h4;
        243: lsb=4'h5;
        244: lsb=4'h0;
        245: lsb=4'h0;
        246: lsb=4'h1;
        247: lsb=4'h2;
        248: lsb=4'h3;
        249: lsb=4'h3;
        250: lsb=4'h4;
        251: lsb=4'h5;
        252: lsb=4'h6;
        253: lsb=4'h7;
        254: lsb=4'hC;
        255: lsb=4'hD;
    endcase

endmodule
