module bit_adder
  (input  a,
   input  b,
   input  ci,
   output s,
   output co);
  wire n1844_o;
  wire n1845_o;
  wire n1846_o;
  wire n1847_o;
  wire n1848_o;
  wire n1849_o;
  wire n1850_o;
  wire n1851_o;
  wire n1852_o;
  wire n1853_o;
  wire n1854_o;
  wire n1855_o;
  wire n1856_o;
  wire n1857_o;
  wire n1858_o;
  wire n1859_o;
  wire n1860_o;
  wire n1861_o;
  wire n1862_o;
  wire n1863_o;
  wire n1864_o;
  wire n1865_o;
  wire n1866_o;
  wire n1867_o;
  wire n1868_o;
  wire n1869_o;
  wire n1870_o;
  wire n1871_o;
  wire n1872_o;
  wire n1873_o;
  wire n1874_o;
  assign s = n1860_o;
  assign co = n1874_o;
  /* AddSubBCD.vhd:21:15  */
  assign n1844_o = ~a;
  /* AddSubBCD.vhd:21:25  */
  assign n1845_o = ~b;
  /* AddSubBCD.vhd:21:21  */
  assign n1846_o = n1844_o & n1845_o;
  /* AddSubBCD.vhd:21:31  */
  assign n1847_o = n1846_o & ci;
  /* AddSubBCD.vhd:22:20  */
  assign n1848_o = ~a;
  /* AddSubBCD.vhd:22:26  */
  assign n1849_o = n1848_o & b;
  /* AddSubBCD.vhd:22:40  */
  assign n1850_o = ~ci;
  /* AddSubBCD.vhd:22:36  */
  assign n1851_o = n1849_o & n1850_o;
  /* AddSubBCD.vhd:21:43  */
  assign n1852_o = n1847_o | n1851_o;
  /* AddSubBCD.vhd:23:30  */
  assign n1853_o = ~b;
  /* AddSubBCD.vhd:23:26  */
  assign n1854_o = a & n1853_o;
  /* AddSubBCD.vhd:23:40  */
  assign n1855_o = ~ci;
  /* AddSubBCD.vhd:23:36  */
  assign n1856_o = n1854_o & n1855_o;
  /* AddSubBCD.vhd:22:48  */
  assign n1857_o = n1852_o | n1856_o;
  /* AddSubBCD.vhd:24:26  */
  assign n1858_o = a & b;
  /* AddSubBCD.vhd:24:36  */
  assign n1859_o = n1858_o & ci;
  /* AddSubBCD.vhd:23:48  */
  assign n1860_o = n1857_o | n1859_o;
  /* AddSubBCD.vhd:26:16  */
  assign n1861_o = ~a;
  /* AddSubBCD.vhd:26:22  */
  assign n1862_o = n1861_o & b;
  /* AddSubBCD.vhd:26:32  */
  assign n1863_o = n1862_o & ci;
  /* AddSubBCD.vhd:27:36  */
  assign n1864_o = ~b;
  /* AddSubBCD.vhd:27:32  */
  assign n1865_o = a & n1864_o;
  /* AddSubBCD.vhd:27:42  */
  assign n1866_o = n1865_o & ci;
  /* AddSubBCD.vhd:26:44  */
  assign n1867_o = n1863_o | n1866_o;
  /* AddSubBCD.vhd:28:32  */
  assign n1868_o = a & b;
  /* AddSubBCD.vhd:28:46  */
  assign n1869_o = ~ci;
  /* AddSubBCD.vhd:28:42  */
  assign n1870_o = n1868_o & n1869_o;
  /* AddSubBCD.vhd:27:54  */
  assign n1871_o = n1867_o | n1870_o;
  /* AddSubBCD.vhd:29:32  */
  assign n1872_o = a & b;
  /* AddSubBCD.vhd:29:42  */
  assign n1873_o = n1872_o & ci;
  /* AddSubBCD.vhd:28:54  */
  assign n1874_o = n1871_o | n1873_o;
endmodule

module adder4
  (input  [3:0] a,
   input  [3:0] b,
   input  ci,
   output [3:0] s,
   output co);
  wire co0;
  wire co1;
  wire co2;
  wire n1809_o;
  wire n1810_o;
  wire b_add0_n1811;
  wire b_add0_n1812;
  wire b_add0_s;
  wire b_add0_co;
  wire n1817_o;
  wire n1818_o;
  wire b_add1_n1819;
  wire b_add1_n1820;
  wire b_add1_s;
  wire b_add1_co;
  wire n1825_o;
  wire n1826_o;
  wire b_add2_n1827;
  wire b_add2_n1828;
  wire b_add2_s;
  wire b_add2_co;
  wire n1833_o;
  wire n1834_o;
  wire b_add3_n1835;
  wire b_add3_n1836;
  wire b_add3_s;
  wire b_add3_co;
  wire [3:0] n1841_o;
  assign s = n1841_o;
  assign co = b_add3_n1836;
  /* AddSubBCD.vhd:63:16  */
  assign co0 = b_add0_n1812; // (signal)
  /* AddSubBCD.vhd:63:21  */
  assign co1 = b_add1_n1820; // (signal)
  /* AddSubBCD.vhd:63:26  */
  assign co2 = b_add2_n1828; // (signal)
  /* AddSubBCD.vhd:67:38  */
  assign n1809_o = a[0];
  /* AddSubBCD.vhd:67:44  */
  assign n1810_o = b[0];
  /* AddSubBCD.vhd:67:54  */
  assign b_add0_n1811 = b_add0_s; // (signal)
  /* AddSubBCD.vhd:67:60  */
  assign b_add0_n1812 = b_add0_co; // (signal)
  /* AddSubBCD.vhd:67:9  */
  bit_adder b_add0 (
    .a(n1809_o),
    .b(n1810_o),
    .ci(ci),
    .s(b_add0_s),
    .co(b_add0_co));
  /* AddSubBCD.vhd:68:38  */
  assign n1817_o = a[1];
  /* AddSubBCD.vhd:68:44  */
  assign n1818_o = b[1];
  /* AddSubBCD.vhd:68:54  */
  assign b_add1_n1819 = b_add1_s; // (signal)
  /* AddSubBCD.vhd:68:60  */
  assign b_add1_n1820 = b_add1_co; // (signal)
  /* AddSubBCD.vhd:68:9  */
  bit_adder b_add1 (
    .a(n1817_o),
    .b(n1818_o),
    .ci(co0),
    .s(b_add1_s),
    .co(b_add1_co));
  /* AddSubBCD.vhd:69:38  */
  assign n1825_o = a[2];
  /* AddSubBCD.vhd:69:44  */
  assign n1826_o = b[2];
  /* AddSubBCD.vhd:69:54  */
  assign b_add2_n1827 = b_add2_s; // (signal)
  /* AddSubBCD.vhd:69:60  */
  assign b_add2_n1828 = b_add2_co; // (signal)
  /* AddSubBCD.vhd:69:9  */
  bit_adder b_add2 (
    .a(n1825_o),
    .b(n1826_o),
    .ci(co1),
    .s(b_add2_s),
    .co(b_add2_co));
  /* AddSubBCD.vhd:70:38  */
  assign n1833_o = a[3];
  /* AddSubBCD.vhd:70:44  */
  assign n1834_o = b[3];
  /* AddSubBCD.vhd:70:54  */
  assign b_add3_n1835 = b_add3_s; // (signal)
  /* AddSubBCD.vhd:70:60  */
  assign b_add3_n1836 = b_add3_co; // (signal)
  /* AddSubBCD.vhd:70:9  */
  bit_adder b_add3 (
    .a(n1833_o),
    .b(n1834_o),
    .ci(co2),
    .s(b_add3_s),
    .co(b_add3_co));
  assign n1841_o = {b_add3_n1835, b_add2_n1827, b_add1_n1819, b_add0_n1811};
endmodule

module bcdadder
  (input  [3:0] a,
   input  [3:0] b,
   input  ci,
   input  add,
   input  bcd,
   output [3:0] s,
   output co,
   output vo);
  wire [3:0] b2;
  wire [3:0] bin_s;
  wire bin_co;
  wire [3:0] bcd_b;
  wire bcd_co;
  wire ci2;
  wire n1764_o;
  wire n1765_o;
  wire n1766_o;
  wire n1767_o;
  wire [3:0] n1768_o;
  wire [3:0] n1769_o;
  wire [3:0] bin_adder_s;
  wire bin_adder_co;
  wire n1772_o;
  wire n1773_o;
  wire n1774_o;
  wire n1775_o;
  wire n1776_o;
  wire n1777_o;
  wire n1778_o;
  wire n1779_o;
  wire n1780_o;
  wire n1781_o;
  wire n1782_o;
  wire n1783_o;
  wire n1784_o;
  wire n1785_o;
  wire [1:0] n1786_o;
  wire n1787_o;
  wire n1788_o;
  wire n1789_o;
  wire [2:0] n1790_o;
  wire n1791_o;
  wire [3:0] n1792_o;
  wire n1793_o;
  wire [3:0] bcd_corr_adder_s;
  wire bcd_corr_adder_co;
  wire n1795_o;
  wire n1796_o;
  wire n1797_o;
  wire n1798_o;
  wire n1799_o;
  wire n1800_o;
  wire n1801_o;
  wire n1802_o;
  wire n1803_o;
  wire n1804_o;
  wire n1805_o;
  wire n1806_o;
  assign s = bcd_corr_adder_s;
  assign co = n1796_o;
  assign vo = n1806_o;
  /* AddSubBCD.vhd:98:16  */
  assign b2 = n1769_o; // (signal)
  /* AddSubBCD.vhd:99:16  */
  assign bin_s = bin_adder_s; // (signal)
  /* AddSubBCD.vhd:100:16  */
  assign bin_co = bin_adder_co; // (signal)
  /* AddSubBCD.vhd:101:16  */
  assign bcd_b = n1792_o; // (signal)
  /* AddSubBCD.vhd:102:16  */
  assign bcd_co = n1781_o; // (signal)
  /* AddSubBCD.vhd:104:16  */
  assign ci2 = n1793_o; // (signal)
  /* AddSubBCD.vhd:108:36  */
  assign n1764_o = ~add;
  /* AddSubBCD.vhd:108:36  */
  assign n1765_o = ~add;
  /* AddSubBCD.vhd:108:36  */
  assign n1766_o = ~add;
  /* AddSubBCD.vhd:108:36  */
  assign n1767_o = ~add;
  assign n1768_o = {n1767_o, n1766_o, n1765_o, n1764_o};
  /* AddSubBCD.vhd:108:17  */
  assign n1769_o = b ^ n1768_o;
  /* AddSubBCD.vhd:110:9  */
  adder4 bin_adder (
    .a(a),
    .b(b2),
    .ci(ci),
    .s(bin_adder_s),
    .co(bin_adder_co));
  /* AddSubBCD.vhd:119:25  */
  assign n1772_o = bin_s[3];
  /* AddSubBCD.vhd:119:38  */
  assign n1773_o = bin_s[2];
  /* AddSubBCD.vhd:119:29  */
  assign n1774_o = n1772_o & n1773_o;
  /* AddSubBCD.vhd:119:52  */
  assign n1775_o = bin_s[3];
  /* AddSubBCD.vhd:119:65  */
  assign n1776_o = bin_s[1];
  /* AddSubBCD.vhd:119:56  */
  assign n1777_o = n1775_o & n1776_o;
  /* AddSubBCD.vhd:119:43  */
  assign n1778_o = n1774_o | n1777_o;
  /* AddSubBCD.vhd:119:85  */
  assign n1779_o = ~add;
  /* AddSubBCD.vhd:119:81  */
  assign n1780_o = bin_co ^ n1779_o;
  /* AddSubBCD.vhd:119:70  */
  assign n1781_o = n1778_o | n1780_o;
  /* AddSubBCD.vhd:120:18  */
  assign n1782_o = ~add;
  /* AddSubBCD.vhd:120:37  */
  assign n1783_o = bcd_co & bcd;
  /* AddSubBCD.vhd:120:50  */
  assign n1784_o = ~add;
  /* AddSubBCD.vhd:120:46  */
  assign n1785_o = n1783_o ^ n1784_o;
  /* AddSubBCD.vhd:120:26  */
  assign n1786_o = {n1782_o, n1785_o};
  /* AddSubBCD.vhd:120:70  */
  assign n1787_o = bcd_co & bcd;
  /* AddSubBCD.vhd:120:83  */
  assign n1788_o = ~add;
  /* AddSubBCD.vhd:120:79  */
  assign n1789_o = n1787_o ^ n1788_o;
  /* AddSubBCD.vhd:120:59  */
  assign n1790_o = {n1786_o, n1789_o};
  /* AddSubBCD.vhd:120:94  */
  assign n1791_o = ~add;
  /* AddSubBCD.vhd:120:92  */
  assign n1792_o = {n1790_o, n1791_o};
  /* AddSubBCD.vhd:122:16  */
  assign n1793_o = ~add;
  /* AddSubBCD.vhd:123:9  */
  adder4 bcd_corr_adder (
    .a(bin_s),
    .b(bcd_b),
    .ci(ci2),
    .s(bcd_corr_adder_s),
    .co());
  /* AddSubBCD.vhd:131:31  */
  assign n1795_o = ~bcd;
  /* AddSubBCD.vhd:131:22  */
  assign n1796_o = n1795_o ? bin_co : n1798_o;
  /* AddSubBCD.vhd:131:53  */
  assign n1797_o = ~add;
  /* AddSubBCD.vhd:131:49  */
  assign n1798_o = bcd_co ^ n1797_o;
  /* AddSubBCD.vhd:132:22  */
  assign n1799_o = a[3];
  /* AddSubBCD.vhd:132:32  */
  assign n1800_o = b2[3];
  /* AddSubBCD.vhd:132:26  */
  assign n1801_o = n1799_o ^ n1800_o;
  /* AddSubBCD.vhd:132:16  */
  assign n1802_o = ~n1801_o;
  /* AddSubBCD.vhd:132:44  */
  assign n1803_o = a[3];
  /* AddSubBCD.vhd:132:57  */
  assign n1804_o = bin_s[3];
  /* AddSubBCD.vhd:132:48  */
  assign n1805_o = n1803_o ^ n1804_o;
  /* AddSubBCD.vhd:132:38  */
  assign n1806_o = n1802_o & n1805_o;
endmodule

module addsubbcd
  (input  [7:0] a,
   input  [7:0] b,
   input  ci,
   input  add,
   input  bcd,
   output [7:0] s,
   output co,
   output vo);
  wire vo1;
  wire co0;
  wire co1;
  wire [3:0] add0_s;
  wire add0_co;
  wire add0_vo;
  wire [3:0] n1751_o;
  wire [3:0] n1752_o;
  wire [3:0] add1_s;
  wire add1_co;
  wire add1_vo;
  wire [3:0] n1755_o;
  wire [3:0] n1756_o;
  wire [7:0] n1760_o;
  assign s = n1760_o;
  assign co = co1;
  assign vo = vo1;
  /* AddSubBCD.vhd:157:16  */
  assign vo1 = add1_vo; // (signal)
  /* AddSubBCD.vhd:158:16  */
  assign co0 = add0_co; // (signal)
  /* AddSubBCD.vhd:158:21  */
  assign co1 = add1_co; // (signal)
  /* AddSubBCD.vhd:162:9  */
  bcdadder add0 (
    .a(n1751_o),
    .b(n1752_o),
    .ci(ci),
    .add(add),
    .bcd(bcd),
    .s(add0_s),
    .co(add0_co),
    .vo());
  /* AddSubBCD.vhd:164:23  */
  assign n1751_o = a[3:0];
  /* AddSubBCD.vhd:165:23  */
  assign n1752_o = b[3:0];
  /* AddSubBCD.vhd:175:9  */
  bcdadder add1 (
    .a(n1755_o),
    .b(n1756_o),
    .ci(co0),
    .add(add),
    .bcd(bcd),
    .s(add1_s),
    .co(add1_co),
    .vo(add1_vo));
  /* AddSubBCD.vhd:177:23  */
  assign n1755_o = a[7:4];
  /* AddSubBCD.vhd:178:23  */
  assign n1756_o = b[7:4];
  assign n1760_o = {add1_s, add0_s};
endmodule

module huc6280_ag
  (input  clk,
   input  rst_n,
   input  ce,
   input  [2:0] pc_ctrl,
   input  [5:0] addr_ctrl,
   input  got_int,
   input  [7:0] di,
   input  [7:0] x,
   input  [7:0] y,
   input  [7:0] dr,
   output [15:0] pc,
   output [15:0] aa);
  wire [7:0] aal;
  wire [7:0] aah;
  wire savedcarry;
  wire [8:0] newaal;
  wire [7:0] newaah;
  wire [15:0] pcr;
  wire [15:0] nextpc;
  wire [15:0] newpcwithoffset;
  wire n1612_o;
  wire n1613_o;
  wire n1614_o;
  wire n1615_o;
  wire n1616_o;
  wire n1617_o;
  wire n1618_o;
  wire n1619_o;
  wire [3:0] n1620_o;
  wire [3:0] n1621_o;
  wire [7:0] n1622_o;
  wire [15:0] n1623_o;
  wire [15:0] n1624_o;
  wire n1628_o;
  wire n1629_o;
  wire [15:0] n1631_o;
  wire [15:0] n1632_o;
  wire n1634_o;
  wire [7:0] n1635_o;
  wire [15:0] n1636_o;
  wire n1638_o;
  wire [7:0] n1639_o;
  wire [15:0] n1640_o;
  wire n1642_o;
  wire n1644_o;
  wire [15:0] n1645_o;
  wire n1647_o;
  wire [5:0] n1648_o;
  reg [15:0] n1649_o;
  wire n1650_o;
  wire [2:0] n1659_o;
  wire [8:0] n1661_o;
  wire n1663_o;
  wire [8:0] n1665_o;
  wire n1667_o;
  wire [8:0] n1669_o;
  wire [8:0] n1671_o;
  wire n1673_o;
  wire [8:0] n1675_o;
  wire [8:0] n1677_o;
  wire [8:0] n1678_o;
  wire n1680_o;
  wire [8:0] n1682_o;
  wire [8:0] n1684_o;
  wire [8:0] n1685_o;
  wire n1687_o;
  wire [8:0] n1689_o;
  wire n1691_o;
  wire [8:0] n1693_o;
  wire [8:0] n1695_o;
  wire [8:0] n1696_o;
  wire n1698_o;
  wire [8:0] n1700_o;
  wire [6:0] n1701_o;
  reg [8:0] n1702_o;
  wire [2:0] n1703_o;
  wire n1705_o;
  wire n1707_o;
  wire [7:0] n1709_o;
  wire n1711_o;
  wire [7:0] n1713_o;
  wire [7:0] n1714_o;
  wire n1716_o;
  wire [3:0] n1717_o;
  reg [7:0] n1718_o;
  wire n1722_o;
  wire [7:0] n1724_o;
  wire n1725_o;
  wire [15:0] n1739_o;
  wire [7:0] n1740_o;
  reg [7:0] n1741_q;
  wire [7:0] n1742_o;
  reg [7:0] n1743_q;
  wire n1744_o;
  reg n1745_q;
  wire [15:0] n1746_o;
  reg [15:0] n1747_q;
  assign pc = pcr;
  assign aa = n1739_o;
  /* HUC6280_AG.vhd:26:16  */
  assign aal = n1741_q; // (signal)
  /* HUC6280_AG.vhd:26:21  */
  assign aah = n1743_q; // (signal)
  /* HUC6280_AG.vhd:27:16  */
  assign savedcarry = n1745_q; // (signal)
  /* HUC6280_AG.vhd:29:16  */
  assign newaal = n1702_o; // (signal)
  /* HUC6280_AG.vhd:117:46  */
  assign newaah = n1718_o; // (signal)
  /* HUC6280_AG.vhd:32:16  */
  assign pcr = n1747_q; // (signal)
  /* HUC6280_AG.vhd:33:16  */
  assign nextpc = n1649_o; // (signal)
  /* HUC6280_AG.vhd:33:24  */
  assign newpcwithoffset = n1624_o; // (signal)
  /* HUC6280_AG.vhd:37:88  */
  assign n1612_o = aal[7];
  /* HUC6280_AG.vhd:37:88  */
  assign n1613_o = aal[7];
  /* HUC6280_AG.vhd:37:88  */
  assign n1614_o = aal[7];
  /* HUC6280_AG.vhd:37:88  */
  assign n1615_o = aal[7];
  /* HUC6280_AG.vhd:37:88  */
  assign n1616_o = aal[7];
  /* HUC6280_AG.vhd:37:88  */
  assign n1617_o = aal[7];
  /* HUC6280_AG.vhd:37:88  */
  assign n1618_o = aal[7];
  /* HUC6280_AG.vhd:37:88  */
  assign n1619_o = aal[7];
  assign n1620_o = {n1619_o, n1618_o, n1617_o, n1616_o};
  assign n1621_o = {n1615_o, n1614_o, n1613_o, n1612_o};
  assign n1622_o = {n1620_o, n1621_o};
  /* HUC6280_AG.vhd:37:93  */
  assign n1623_o = {n1622_o, aal};
  /* HUC6280_AG.vhd:37:59  */
  assign n1624_o = pcr + n1623_o;
  /* HUC6280_AG.vhd:42:25  */
  assign n1628_o = pc_ctrl == 3'b000;
  /* HUC6280_AG.vhd:45:44  */
  assign n1629_o = ~got_int;
  /* HUC6280_AG.vhd:46:82  */
  assign n1631_o = pcr + 16'b0000000000000001;
  /* HUC6280_AG.vhd:45:33  */
  assign n1632_o = n1629_o ? n1631_o : pcr;
  /* HUC6280_AG.vhd:44:25  */
  assign n1634_o = pc_ctrl == 3'b001;
  /* HUC6280_AG.vhd:51:46  */
  assign n1635_o = pcr[15:8];
  /* HUC6280_AG.vhd:51:60  */
  assign n1636_o = {n1635_o, di};
  /* HUC6280_AG.vhd:50:25  */
  assign n1638_o = pc_ctrl == 3'b010;
  /* HUC6280_AG.vhd:53:51  */
  assign n1639_o = pcr[7:0];
  /* HUC6280_AG.vhd:53:46  */
  assign n1640_o = {di, n1639_o};
  /* HUC6280_AG.vhd:52:25  */
  assign n1642_o = pc_ctrl == 3'b011;
  /* HUC6280_AG.vhd:54:25  */
  assign n1644_o = pc_ctrl == 3'b100;
  /* HUC6280_AG.vhd:57:47  */
  assign n1645_o = {aah, aal};
  /* HUC6280_AG.vhd:56:25  */
  assign n1647_o = pc_ctrl == 3'b110;
  assign n1648_o = {n1647_o, n1644_o, n1642_o, n1638_o, n1634_o, n1628_o};
  /* HUC6280_AG.vhd:41:17  */
  always @*
    case (n1648_o)
      6'b100000: n1649_o = n1645_o;
      6'b010000: n1649_o = newpcwithoffset;
      6'b001000: n1649_o = n1640_o;
      6'b000100: n1649_o = n1636_o;
      6'b000010: n1649_o = n1632_o;
      6'b000001: n1649_o = pcr;
      default: n1649_o = pcr;
    endcase
  /* HUC6280_AG.vhd:62:26  */
  assign n1650_o = ~rst_n;
  /* HUC6280_AG.vhd:73:31  */
  assign n1659_o = addr_ctrl[5:3];
  /* HUC6280_AG.vhd:75:47  */
  assign n1661_o = {1'b0, aal};
  /* HUC6280_AG.vhd:74:25  */
  assign n1663_o = n1659_o == 3'b000;
  /* HUC6280_AG.vhd:77:47  */
  assign n1665_o = {1'b0, di};
  /* HUC6280_AG.vhd:76:25  */
  assign n1667_o = n1659_o == 3'b001;
  /* HUC6280_AG.vhd:79:73  */
  assign n1669_o = {1'b0, aal};
  /* HUC6280_AG.vhd:79:80  */
  assign n1671_o = n1669_o + 9'b000000001;
  /* HUC6280_AG.vhd:78:25  */
  assign n1673_o = n1659_o == 3'b010;
  /* HUC6280_AG.vhd:81:73  */
  assign n1675_o = {1'b0, aal};
  /* HUC6280_AG.vhd:81:95  */
  assign n1677_o = {1'b0, x};
  /* HUC6280_AG.vhd:81:80  */
  assign n1678_o = n1675_o + n1677_o;
  /* HUC6280_AG.vhd:80:25  */
  assign n1680_o = n1659_o == 3'b011;
  /* HUC6280_AG.vhd:83:73  */
  assign n1682_o = {1'b0, aal};
  /* HUC6280_AG.vhd:83:95  */
  assign n1684_o = {1'b0, y};
  /* HUC6280_AG.vhd:83:80  */
  assign n1685_o = n1682_o + n1684_o;
  /* HUC6280_AG.vhd:82:25  */
  assign n1687_o = n1659_o == 3'b100;
  /* HUC6280_AG.vhd:85:47  */
  assign n1689_o = {1'b0, dr};
  /* HUC6280_AG.vhd:84:25  */
  assign n1691_o = n1659_o == 3'b101;
  /* HUC6280_AG.vhd:87:73  */
  assign n1693_o = {1'b0, dr};
  /* HUC6280_AG.vhd:87:94  */
  assign n1695_o = {1'b0, y};
  /* HUC6280_AG.vhd:87:79  */
  assign n1696_o = n1693_o + n1695_o;
  /* HUC6280_AG.vhd:86:25  */
  assign n1698_o = n1659_o == 3'b110;
  /* HUC6280_AG.vhd:89:47  */
  assign n1700_o = {1'b0, x};
  assign n1701_o = {n1698_o, n1691_o, n1687_o, n1680_o, n1673_o, n1667_o, n1663_o};
  /* HUC6280_AG.vhd:73:17  */
  always @*
    case (n1701_o)
      7'b1000000: n1702_o = n1696_o;
      7'b0100000: n1702_o = n1689_o;
      7'b0010000: n1702_o = n1685_o;
      7'b0001000: n1702_o = n1678_o;
      7'b0000100: n1702_o = n1671_o;
      7'b0000010: n1702_o = n1665_o;
      7'b0000001: n1702_o = n1661_o;
      default: n1702_o = n1700_o;
    endcase
  /* HUC6280_AG.vhd:92:31  */
  assign n1703_o = addr_ctrl[2:0];
  /* HUC6280_AG.vhd:93:25  */
  assign n1705_o = n1703_o == 3'b000;
  /* HUC6280_AG.vhd:95:25  */
  assign n1707_o = n1703_o == 3'b001;
  /* HUC6280_AG.vhd:98:74  */
  assign n1709_o = aah + 8'b00000001;
  /* HUC6280_AG.vhd:97:25  */
  assign n1711_o = n1703_o == 3'b010;
  /* HUC6280_AG.vhd:100:86  */
  assign n1713_o = {7'b0000000, savedcarry};
  /* HUC6280_AG.vhd:100:74  */
  assign n1714_o = aah + n1713_o;
  /* HUC6280_AG.vhd:99:25  */
  assign n1716_o = n1703_o == 3'b011;
  assign n1717_o = {n1716_o, n1711_o, n1707_o, n1705_o};
  /* HUC6280_AG.vhd:92:17  */
  always @*
    case (n1717_o)
      4'b1000: n1718_o = n1714_o;
      4'b0100: n1718_o = n1709_o;
      4'b0010: n1718_o = di;
      4'b0001: n1718_o = aah;
      default: n1718_o = aah;
    endcase
  /* HUC6280_AG.vhd:109:26  */
  assign n1722_o = ~rst_n;
  /* HUC6280_AG.vhd:115:46  */
  assign n1724_o = newaal[7:0];
  /* HUC6280_AG.vhd:116:53  */
  assign n1725_o = newaal[8];
  /* HUC6280_AG.vhd:122:19  */
  assign n1739_o = {aah, aal};
  /* HUC6280_AG.vhd:113:17  */
  assign n1740_o = ce ? n1724_o : aal;
  /* HUC6280_AG.vhd:113:17  */
  always @(posedge clk or posedge n1722_o)
    if (n1722_o)
      n1741_q <= 8'b00000000;
    else
      n1741_q <= n1740_o;
  /* HUC6280_AG.vhd:113:17  */
  assign n1742_o = ce ? newaah : aah;
  /* HUC6280_AG.vhd:113:17  */
  always @(posedge clk or posedge n1722_o)
    if (n1722_o)
      n1743_q <= 8'b00000000;
    else
      n1743_q <= n1742_o;
  /* HUC6280_AG.vhd:113:17  */
  assign n1744_o = ce ? n1725_o : savedcarry;
  /* HUC6280_AG.vhd:113:17  */
  always @(posedge clk or posedge n1722_o)
    if (n1722_o)
      n1745_q <= 1'b0;
    else
      n1745_q <= n1744_o;
  /* HUC6280_AG.vhd:64:17  */
  assign n1746_o = ce ? nextpc : pcr;
  /* HUC6280_AG.vhd:64:17  */
  always @(posedge clk or posedge n1650_o)
    if (n1650_o)
      n1747_q <= 16'b0000000000000000;
    else
      n1747_q <= n1746_o;
endmodule

module alu
  (input  clk,
   input  en,
   input  [7:0] l,
   input  [7:0] r,
   input  [2:0] ctrl_fstop,
   input  [2:0] ctrl_secop,
   input  ctrl_fc,
   input  bcd,
   input  ci,
   input  vi,
   input  ni,
   output co,
   output vo,
   output no,
   output zo,
   output [7:0] res);
  wire [6:0] n1470_o;
  wire [7:0] intl;
  wire [7:0] intr;
  wire cr;
  wire addin;
  wire bcdin;
  wire ciin;
  wire savedc;
  wire [7:0] adds;
  wire addco;
  wire addvo;
  wire [7:0] result;
  wire [2:0] n1478_o;
  wire n1479_o;
  wire [6:0] n1480_o;
  wire [7:0] n1482_o;
  wire n1484_o;
  wire n1485_o;
  wire [6:0] n1486_o;
  wire [7:0] n1487_o;
  wire n1489_o;
  wire n1490_o;
  wire [6:0] n1491_o;
  wire [7:0] n1493_o;
  wire n1495_o;
  wire n1496_o;
  wire [6:0] n1497_o;
  wire [7:0] n1498_o;
  wire n1500_o;
  wire n1501_o;
  wire n1502_o;
  wire n1503_o;
  wire n1504_o;
  wire n1506_o;
  wire n1508_o;
  wire n1509_o;
  wire n1511_o;
  wire n1513_o;
  wire [7:0] n1514_o;
  reg [7:0] n1515_o;
  reg [7:0] n1522_o;
  reg n1523_o;
  reg n1525_o;
  wire n1528_o;
  wire n1529_o;
  wire n1530_o;
  wire n1531_o;
  wire n1532_o;
  wire [7:0] addsub_s;
  wire addsub_co;
  wire addsub_vo;
  wire [2:0] n1544_o;
  wire [7:0] n1545_o;
  wire n1547_o;
  wire [7:0] n1548_o;
  wire n1550_o;
  wire [7:0] n1551_o;
  wire n1553_o;
  wire n1555_o;
  wire n1557_o;
  wire n1558_o;
  wire n1560_o;
  wire n1561_o;
  wire n1563_o;
  wire n1564_o;
  wire n1565_o;
  wire [7:0] n1566_o;
  wire [7:0] n1567_o;
  wire [7:0] n1568_o;
  wire [7:0] n1569_o;
  wire n1571_o;
  wire [5:0] n1572_o;
  reg n1573_o;
  reg [7:0] n1574_o;
  wire n1578_o;
  wire [2:0] n1579_o;
  wire n1580_o;
  wire n1581_o;
  wire n1582_o;
  wire n1583_o;
  wire n1584_o;
  wire n1586_o;
  wire n1587_o;
  wire n1588_o;
  wire n1590_o;
  wire n1591_o;
  wire n1592_o;
  wire n1594_o;
  wire n1595_o;
  wire n1596_o;
  wire n1598_o;
  wire [3:0] n1599_o;
  reg n1600_o;
  reg n1601_o;
  wire n1605_o;
  wire n1606_o;
  wire n1608_o;
  reg n1609_q;
  assign co = n1573_o;
  assign vo = n1600_o;
  assign no = n1601_o;
  assign zo = n1606_o;
  assign res = result;
  /* HUC6280_MC.vhd:6978:17  */
  assign n1470_o = {ctrl_fc, ctrl_secop, ctrl_fstop};
  /* HUC6280_ALU.vhd:28:16  */
  assign intl = n1515_o; // (signal)
  /* HUC6280_ALU.vhd:29:16  */
  assign intr = n1522_o; // (signal)
  /* HUC6280_ALU.vhd:30:16  */
  assign cr = n1523_o; // (signal)
  /* HUC6280_ALU.vhd:31:16  */
  assign addin = n1532_o; // (signal)
  /* HUC6280_ALU.vhd:32:16  */
  assign bcdin = n1525_o; // (signal)
  /* HUC6280_ALU.vhd:33:16  */
  assign ciin = n1530_o; // (signal)
  /* HUC6280_ALU.vhd:34:16  */
  assign savedc = n1609_q; // (signal)
  /* HUC6280_ALU.vhd:36:16  */
  assign adds = addsub_s; // (signal)
  /* HUC6280_ALU.vhd:37:16  */
  assign addco = addsub_co; // (signal)
  /* HUC6280_ALU.vhd:38:16  */
  assign addvo = addsub_vo; // (signal)
  /* HUC6280_ALU.vhd:39:16  */
  assign result = n1574_o; // (signal)
  /* HUC6280_ALU.vhd:47:27  */
  assign n1478_o = n1470_o[2:0];
  /* HUC6280_ALU.vhd:49:40  */
  assign n1479_o = l[7];
  /* HUC6280_ALU.vhd:50:42  */
  assign n1480_o = l[6:0];
  /* HUC6280_ALU.vhd:50:55  */
  assign n1482_o = {n1480_o, 1'b0};
  /* HUC6280_ALU.vhd:48:25  */
  assign n1484_o = n1478_o == 3'b000;
  /* HUC6280_ALU.vhd:53:40  */
  assign n1485_o = l[7];
  /* HUC6280_ALU.vhd:54:42  */
  assign n1486_o = l[6:0];
  /* HUC6280_ALU.vhd:54:55  */
  assign n1487_o = {n1486_o, ci};
  /* HUC6280_ALU.vhd:52:25  */
  assign n1489_o = n1478_o == 3'b001;
  /* HUC6280_ALU.vhd:57:40  */
  assign n1490_o = l[0];
  /* HUC6280_ALU.vhd:58:48  */
  assign n1491_o = l[7:1];
  /* HUC6280_ALU.vhd:58:45  */
  assign n1493_o = {1'b0, n1491_o};
  /* HUC6280_ALU.vhd:56:25  */
  assign n1495_o = n1478_o == 3'b010;
  /* HUC6280_ALU.vhd:61:40  */
  assign n1496_o = l[0];
  /* HUC6280_ALU.vhd:62:47  */
  assign n1497_o = l[7:1];
  /* HUC6280_ALU.vhd:62:44  */
  assign n1498_o = {ci, n1497_o};
  /* HUC6280_ALU.vhd:60:25  */
  assign n1500_o = n1478_o == 3'b011;
  /* HUC6280_ALU.vhd:67:60  */
  assign n1501_o = n1470_o[4];
  /* HUC6280_ALU.vhd:67:46  */
  assign n1502_o = bcd & n1501_o;
  /* HUC6280_ALU.vhd:67:78  */
  assign n1503_o = n1470_o[3];
  /* HUC6280_ALU.vhd:67:64  */
  assign n1504_o = n1502_o & n1503_o;
  /* HUC6280_ALU.vhd:64:25  */
  assign n1506_o = n1478_o == 3'b100;
  /* HUC6280_ALU.vhd:68:25  */
  assign n1508_o = n1478_o == 3'b101;
  /* HUC6280_ALU.vhd:74:49  */
  assign n1509_o = n1470_o[5];
  /* HUC6280_ALU.vhd:71:25  */
  assign n1511_o = n1478_o == 3'b110;
  /* HUC6280_ALU.vhd:75:25  */
  assign n1513_o = n1478_o == 3'b111;
  assign n1514_o = {n1513_o, n1511_o, n1508_o, n1506_o, n1500_o, n1495_o, n1489_o, n1484_o};
  /* HUC6280_ALU.vhd:47:17  */
  always @*
    case (n1514_o)
      8'b10000000: n1515_o = l;
      8'b01000000: n1515_o = l;
      8'b00100000: n1515_o = l;
      8'b00010000: n1515_o = l;
      8'b00001000: n1515_o = n1498_o;
      8'b00000100: n1515_o = n1493_o;
      8'b00000010: n1515_o = n1487_o;
      8'b00000001: n1515_o = n1482_o;
      default: n1515_o = intl;
    endcase
  /* HUC6280_ALU.vhd:47:17  */
  always @*
    case (n1514_o)
      8'b10000000: n1522_o = 8'b00000000;
      8'b01000000: n1522_o = 8'b00000001;
      8'b00100000: n1522_o = r;
      8'b00010000: n1522_o = r;
      8'b00001000: n1522_o = 8'b00000000;
      8'b00000100: n1522_o = 8'b00000000;
      8'b00000010: n1522_o = 8'b00000000;
      8'b00000001: n1522_o = 8'b00000000;
      default: n1522_o = intr;
    endcase
  /* HUC6280_ALU.vhd:47:17  */
  always @*
    case (n1514_o)
      8'b10000000: n1523_o = savedc;
      8'b01000000: n1523_o = n1509_o;
      8'b00100000: n1523_o = ci;
      8'b00010000: n1523_o = ci;
      8'b00001000: n1523_o = n1496_o;
      8'b00000100: n1523_o = n1490_o;
      8'b00000010: n1523_o = n1485_o;
      8'b00000001: n1523_o = n1479_o;
      default: n1523_o = ci;
    endcase
  /* HUC6280_ALU.vhd:47:17  */
  always @*
    case (n1514_o)
      8'b10000000: n1525_o = 1'b0;
      8'b01000000: n1525_o = 1'b0;
      8'b00100000: n1525_o = 1'b0;
      8'b00010000: n1525_o = n1504_o;
      8'b00001000: n1525_o = 1'b0;
      8'b00000100: n1525_o = 1'b0;
      8'b00000010: n1525_o = 1'b0;
      8'b00000001: n1525_o = 1'b0;
      default: n1525_o = 1'b0;
    endcase
  /* HUC6280_ALU.vhd:83:37  */
  assign n1528_o = n1470_o[3];
  /* HUC6280_ALU.vhd:83:23  */
  assign n1529_o = ~n1528_o;
  /* HUC6280_ALU.vhd:83:20  */
  assign n1530_o = cr | n1529_o;
  /* HUC6280_ALU.vhd:84:32  */
  assign n1531_o = n1470_o[5];
  /* HUC6280_ALU.vhd:84:18  */
  assign n1532_o = ~n1531_o;
  /* HUC6280_ALU.vhd:86:9  */
  addsubbcd addsub (
    .a(intl),
    .b(intr),
    .ci(ciin),
    .add(addin),
    .bcd(bcdin),
    .s(addsub_s),
    .co(addsub_co),
    .vo(addsub_vo));
  /* HUC6280_ALU.vhd:109:27  */
  assign n1544_o = n1470_o[5:3];
  /* HUC6280_ALU.vhd:112:48  */
  assign n1545_o = intl | intr;
  /* HUC6280_ALU.vhd:110:25  */
  assign n1547_o = n1544_o == 3'b000;
  /* HUC6280_ALU.vhd:115:48  */
  assign n1548_o = intl & intr;
  /* HUC6280_ALU.vhd:113:25  */
  assign n1550_o = n1544_o == 3'b001;
  /* HUC6280_ALU.vhd:118:48  */
  assign n1551_o = intl ^ intr;
  /* HUC6280_ALU.vhd:116:25  */
  assign n1553_o = n1544_o == 3'b010;
  /* HUC6280_ALU.vhd:119:25  */
  assign n1555_o = n1544_o == 3'b011;
  /* HUC6280_ALU.vhd:119:36  */
  assign n1557_o = n1544_o == 3'b110;
  /* HUC6280_ALU.vhd:119:36  */
  assign n1558_o = n1555_o | n1557_o;
  /* HUC6280_ALU.vhd:119:44  */
  assign n1560_o = n1544_o == 3'b111;
  /* HUC6280_ALU.vhd:119:44  */
  assign n1561_o = n1558_o | n1560_o;
  /* HUC6280_ALU.vhd:122:25  */
  assign n1563_o = n1544_o == 3'b100;
  /* HUC6280_ALU.vhd:127:41  */
  assign n1564_o = n1470_o[6];
  /* HUC6280_ALU.vhd:127:44  */
  assign n1565_o = ~n1564_o;
  /* HUC6280_ALU.vhd:128:61  */
  assign n1566_o = ~intl;
  /* HUC6280_ALU.vhd:128:56  */
  assign n1567_o = intr & n1566_o;
  /* HUC6280_ALU.vhd:130:56  */
  assign n1568_o = intr | intl;
  /* HUC6280_ALU.vhd:127:33  */
  assign n1569_o = n1565_o ? n1567_o : n1568_o;
  /* HUC6280_ALU.vhd:125:25  */
  assign n1571_o = n1544_o == 3'b101;
  assign n1572_o = {n1571_o, n1563_o, n1561_o, n1553_o, n1550_o, n1547_o};
  /* HUC6280_ALU.vhd:109:17  */
  always @*
    case (n1572_o)
      6'b100000: n1573_o = cr;
      6'b010000: n1573_o = cr;
      6'b001000: n1573_o = addco;
      6'b000100: n1573_o = cr;
      6'b000010: n1573_o = cr;
      6'b000001: n1573_o = cr;
      default: n1573_o = n1573_o;
    endcase
  /* HUC6280_ALU.vhd:109:17  */
  always @*
    case (n1572_o)
      6'b100000: n1574_o = n1569_o;
      6'b010000: n1574_o = intl;
      6'b001000: n1574_o = adds;
      6'b000100: n1574_o = n1551_o;
      6'b000010: n1574_o = n1548_o;
      6'b000001: n1574_o = n1545_o;
      default: n1574_o = result;
    endcase
  /* HUC6280_ALU.vhd:139:29  */
  assign n1578_o = result[7];
  /* HUC6280_ALU.vhd:140:27  */
  assign n1579_o = n1470_o[5:3];
  /* HUC6280_ALU.vhd:142:41  */
  assign n1580_o = n1470_o[6];
  /* HUC6280_ALU.vhd:143:51  */
  assign n1581_o = intr[6];
  /* HUC6280_ALU.vhd:144:51  */
  assign n1582_o = intr[7];
  /* HUC6280_ALU.vhd:142:33  */
  assign n1583_o = n1580_o ? n1581_o : vi;
  /* HUC6280_ALU.vhd:142:33  */
  assign n1584_o = n1580_o ? n1582_o : n1578_o;
  /* HUC6280_ALU.vhd:141:25  */
  assign n1586_o = n1579_o == 3'b001;
  /* HUC6280_ALU.vhd:147:42  */
  assign n1587_o = ~bcdin;
  /* HUC6280_ALU.vhd:147:33  */
  assign n1588_o = n1587_o ? addvo : vi;
  /* HUC6280_ALU.vhd:146:25  */
  assign n1590_o = n1579_o == 3'b011;
  /* HUC6280_ALU.vhd:151:43  */
  assign n1591_o = intr[6];
  /* HUC6280_ALU.vhd:152:43  */
  assign n1592_o = intr[7];
  /* HUC6280_ALU.vhd:150:25  */
  assign n1594_o = n1579_o == 3'b101;
  /* HUC6280_ALU.vhd:154:42  */
  assign n1595_o = ~bcdin;
  /* HUC6280_ALU.vhd:154:33  */
  assign n1596_o = n1595_o ? addvo : vi;
  /* HUC6280_ALU.vhd:153:25  */
  assign n1598_o = n1579_o == 3'b111;
  assign n1599_o = {n1598_o, n1594_o, n1590_o, n1586_o};
  /* HUC6280_ALU.vhd:140:17  */
  always @*
    case (n1599_o)
      4'b1000: n1600_o = n1596_o;
      4'b0100: n1600_o = n1591_o;
      4'b0010: n1600_o = n1588_o;
      4'b0001: n1600_o = n1583_o;
      default: n1600_o = vi;
    endcase
  /* HUC6280_ALU.vhd:140:17  */
  always @*
    case (n1599_o)
      4'b1000: n1601_o = n1578_o;
      4'b0100: n1601_o = n1592_o;
      4'b0010: n1601_o = n1578_o;
      4'b0001: n1601_o = n1584_o;
      default: n1601_o = n1578_o;
    endcase
  /* HUC6280_ALU.vhd:162:31  */
  assign n1605_o = result == 8'b00000000;
  /* HUC6280_ALU.vhd:162:19  */
  assign n1606_o = n1605_o ? 1'b1 : 1'b0;
  /* HUC6280_ALU.vhd:100:17  */
  assign n1608_o = en ? addco : savedc;
  /* HUC6280_ALU.vhd:100:17  */
  always @(posedge clk)
    n1609_q <= n1608_o;
endmodule

module huc6280_mc
  (input  clk,
   input  rst_n,
   input  en,
   input  [7:0] ir,
   input  [4:0] state,
   output [1:0] m_state_ctrl,
   output [2:0] m_addr_bus,
   output [1:0] m_load_sdlh,
   output [2:0] m_load_p,
   output [2:0] m_load_t,
   output [5:0] m_addr_ctrl,
   output [2:0] m_load_pc,
   output [2:0] m_load_sp,
   output [2:0] m_axy_ctrl,
   output [3:0] m_alubus_ctrl,
   output [3:0] m_out_bus,
   output m_mem_cycle,
   output [6:0] m_alu_ctrl);
  wire [1:0] n1371_o;
  wire [2:0] n1372_o;
  wire [1:0] n1373_o;
  wire [2:0] n1374_o;
  wire [2:0] n1375_o;
  wire [5:0] n1376_o;
  wire [2:0] n1377_o;
  wire [2:0] n1378_o;
  wire [2:0] n1379_o;
  wire [3:0] n1380_o;
  wire [3:0] n1381_o;
  wire n1382_o;
  wire [6:0] n1383_o;
  wire [41:0] mi;
  wire [6:0] aluflags;
  wire [4:0] n1384_o;
  wire [4:0] n1387_o;
  wire n1394_o;
  wire [2:0] n1396_o;
  wire [10:0] n1397_o;
  wire n1399_o;
  wire [1:0] n1400_o;
  wire n1402_o;
  wire [10:0] n1405_o;
  wire [1:0] n1409_o;
  wire n1411_o;
  wire [10:0] n1414_o;
  wire [1:0] n1418_o;
  wire n1420_o;
  wire [10:0] n1423_o;
  wire [41:0] n1427_o;
  wire [41:0] n1428_o;
  wire [41:0] n1429_o;
  wire [41:0] n1431_o;
  wire [1:0] n1444_o;
  wire [2:0] n1445_o;
  wire [1:0] n1446_o;
  wire [2:0] n1447_o;
  wire [2:0] n1448_o;
  wire [5:0] n1449_o;
  wire [2:0] n1450_o;
  wire [2:0] n1451_o;
  wire [2:0] n1452_o;
  wire [3:0] n1453_o;
  wire [3:0] n1454_o;
  wire n1455_o;
  wire [15:0] n1456_o;
  wire [14:0] n1457_o;
  wire [10:0] n1458_o;
  wire [43:0] n1459_o;
  wire [41:0] n1460_o;
  reg [41:0] n1461_q;
  wire [6:0] n1463_data; // mem_rd
  wire [41:0] n1465_data; // mem_rd
  wire [41:0] n1467_data; // mem_rd
  wire [41:0] n1469_data; // mem_rd
  assign m_state_ctrl = n1371_o;
  assign m_addr_bus = n1372_o;
  assign m_load_sdlh = n1373_o;
  assign m_load_p = n1374_o;
  assign m_load_t = n1375_o;
  assign m_addr_ctrl = n1376_o;
  assign m_load_pc = n1377_o;
  assign m_load_sp = n1378_o;
  assign m_axy_ctrl = n1379_o;
  assign m_alubus_ctrl = n1380_o;
  assign m_out_bus = n1381_o;
  assign m_mem_cycle = n1382_o;
  assign m_alu_ctrl = n1383_o;
  /* HUC6280_CPU.vhd:482:17  */
  assign n1371_o = n1459_o[1:0];
  /* HUC6280_CPU.vhd:472:9  */
  assign n1372_o = n1459_o[4:2];
  assign n1373_o = n1459_o[6:5];
  /* HUC6280_CPU.vhd:460:17  */
  assign n1374_o = n1459_o[9:7];
  /* HUC6280_CPU.vhd:460:17  */
  assign n1375_o = n1459_o[12:10];
  /* HUC6280_CPU.vhd:455:9  */
  assign n1376_o = n1459_o[18:13];
  assign n1377_o = n1459_o[21:19];
  /* HUC6280_CPU.vhd:431:17  */
  assign n1378_o = n1459_o[24:22];
  /* HUC6280_CPU.vhd:427:9  */
  assign n1379_o = n1459_o[27:25];
  assign n1380_o = n1459_o[31:28];
  assign n1381_o = n1459_o[35:32];
  /* HUC6280_CPU.vhd:419:9  */
  assign n1382_o = n1459_o[36];
  assign n1383_o = n1459_o[43:37];
  /* HUC6280_MC.vhd:6966:16  */
  assign mi = n1461_q; // (signal)
  /* HUC6280_MC.vhd:6967:16  */
  assign aluflags = n1463_data; // (signal)
  /* HUC6280_MC.vhd:6971:52  */
  assign n1384_o = mi[36:32];
  /* HUC6280_MC.vhd:6971:29  */
  assign n1387_o = 5'b10001 - n1384_o;
  /* HUC6280_MC.vhd:6976:26  */
  assign n1394_o = ~rst_n;
  /* HUC6280_MC.vhd:6980:56  */
  assign n1396_o = state[2:0];
  /* HUC6280_MC.vhd:6980:50  */
  assign n1397_o = {ir, n1396_o};
  /* HUC6280_MC.vhd:6981:42  */
  assign n1399_o = state == 5'b00000;
  /* HUC6280_MC.vhd:6983:44  */
  assign n1400_o = state[4:3];
  /* HUC6280_MC.vhd:6983:57  */
  assign n1402_o = n1400_o == 2'b00;
  /* HUC6280_MC.vhd:6984:54  */
  assign n1405_o = 11'b11111111111 - n1397_o;
  /* HUC6280_MC.vhd:6985:44  */
  assign n1409_o = state[4:3];
  /* HUC6280_MC.vhd:6985:57  */
  assign n1411_o = n1409_o == 2'b01;
  /* HUC6280_MC.vhd:6986:54  */
  assign n1414_o = 11'b11111111111 - n1397_o;
  /* HUC6280_MC.vhd:6987:44  */
  assign n1418_o = state[4:3];
  /* HUC6280_MC.vhd:6987:57  */
  assign n1420_o = n1418_o == 2'b10;
  /* HUC6280_MC.vhd:6988:54  */
  assign n1423_o = 11'b11111111111 - n1397_o;
  /* HUC6280_MC.vhd:6987:33  */
  assign n1427_o = n1420_o ? n1469_data : mi;
  /* HUC6280_MC.vhd:6985:33  */
  assign n1428_o = n1411_o ? n1467_data : n1427_o;
  /* HUC6280_MC.vhd:6983:33  */
  assign n1429_o = n1402_o ? n1465_data : n1428_o;
  /* HUC6280_MC.vhd:6981:33  */
  assign n1431_o = n1399_o ? 42'b100000000000000000000010000000000000000000 : n1429_o;
  /* HUC6280_MC.vhd:6994:18  */
  assign n1444_o = mi[1:0];
  /* HUC6280_MC.vhd:6995:28  */
  assign n1445_o = mi[4:2];
  /* HUC6280_MC.vhd:6996:28  */
  assign n1446_o = mi[6:5];
  /* HUC6280_MC.vhd:6997:28  */
  assign n1447_o = mi[9:7];
  /* HUC6280_MC.vhd:6998:28  */
  assign n1448_o = mi[12:10];
  /* HUC6280_MC.vhd:6999:28  */
  assign n1449_o = mi[18:13];
  /* HUC6280_MC.vhd:7000:28  */
  assign n1450_o = mi[21:19];
  /* HUC6280_MC.vhd:7001:28  */
  assign n1451_o = mi[24:22];
  /* HUC6280_MC.vhd:7002:28  */
  assign n1452_o = mi[27:25];
  /* HUC6280_MC.vhd:7003:28  */
  assign n1453_o = mi[31:28];
  /* HUC6280_MC.vhd:7004:28  */
  assign n1454_o = mi[40:37];
  /* HUC6280_MC.vhd:7005:28  */
  assign n1455_o = mi[41];
  assign n1456_o = {aluflags, n1455_o, n1454_o, n1453_o};
  assign n1457_o = {n1452_o, n1451_o, n1450_o, n1449_o};
  assign n1458_o = {n1448_o, n1447_o, n1446_o, n1445_o};
  assign n1459_o = {n1456_o, n1457_o, n1458_o, n1444_o};
  /* HUC6280_MC.vhd:6978:17  */
  assign n1460_o = en ? n1431_o : mi;
  /* HUC6280_MC.vhd:6978:17  */
  always @(posedge clk or posedge n1394_o)
    if (n1394_o)
      n1461_q <= 42'b100000000000000000000010000000000000000000;
    else
      n1461_q <= n1460_o;
  /* HUC6280_MC.vhd:14:9  */
  reg [6:0] n1462[17:0] ; // memory
  initial begin
    n1462[17] = 7'b0100100;
    n1462[16] = 7'b0001100;
    n1462[15] = 7'b0000100;
    n1462[14] = 7'b0010100;
    n1462[13] = 7'b0011100;
    n1462[12] = 7'b1111100;
    n1462[11] = 7'b0111110;
    n1462[10] = 7'b0011110;
    n1462[9] = 7'b0100000;
    n1462[8] = 7'b0100010;
    n1462[7] = 7'b0100001;
    n1462[6] = 7'b0100011;
    n1462[5] = 7'b1001100;
    n1462[4] = 7'b0101100;
    n1462[3] = 7'b1101100;
    n1462[2] = 7'b0110100;
    n1462[1] = 7'b0111111;
    n1462[0] = 7'b0011111;
    end
  assign n1463_data = n1462[n1387_o];
  /* HUC6280_MC.vhd:6971:29  */
  /* HUC6280_MC.vhd:6971:28  */
  reg [41:0] n1464[2047:0] ; // memory
  initial begin
    n1464[2047] = 42'b100000000000000000000010000000000000000000;
    n1464[2046] = 42'b100000000000000000000010000000000000000000;
    n1464[2045] = 42'b000000000000000000000000000000000000000000;
    n1464[2044] = 42'b101100000000000000110000000000000000001000;
    n1464[2043] = 42'b101110000000000000110000000000000000001000;
    n1464[2042] = 42'b101010000000000000110000000000000000001000;
    n1464[2041] = 42'b100000000000000000000100000000000100010000;
    n1464[2040] = 42'b100000000000000000000110000000000000010010;
    n1464[2039] = 42'b100000000000000000000010000000000000000000;
    n1464[2038] = 42'b100000000000000000000010010000000000000000;
    n1464[2037] = 42'b000000000000000000000000110000000000000000;
    n1464[2036] = 42'b100000000000000000000000100000000000001100;
    n1464[2035] = 42'b100000000000000000000001010010000000001100;
    n1464[2034] = 42'b000000000000000000000000000000000000000000;
    n1464[2033] = 42'b100000001000010010000000000000000010000110;
    n1464[2032] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2031] = 42'b100000000000000000000010000000000000000000;
    n1464[2030] = 42'b100000000000110100000000000000100000000000;
    n1464[2029] = 42'b000000000001011000000000000000000000000010;
    n1464[2028] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2027] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2026] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2025] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2024] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2023] = 42'b100000000000000000000010000000000000000000;
    n1464[2022] = 42'b100000000000000000000010000000010000000000;
    n1464[2021] = 42'b000000000000000000000000000000000000000000;
    n1464[2020] = 42'b101000000000000000000000000000000000010110;
    n1464[2019] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2018] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2017] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2016] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2015] = 42'b100000000000000000000010000000000000000000;
    n1464[2014] = 42'b100000000000000000000010010000000000000000;
    n1464[2013] = 42'b000000000000000000000000000000000000000000;
    n1464[2012] = 42'b100000111000010000000000000000011010001100;
    n1464[2011] = 42'b000000000000000000000000000000000000000000;
    n1464[2010] = 42'b101000000000000000000000000000000000001110;
    n1464[2009] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2008] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2007] = 42'b100000000000000000000010000000000000000000;
    n1464[2006] = 42'b100000000000000000000010010000000000000000;
    n1464[2005] = 42'b000000000000000000000000000000000000000000;
    n1464[2004] = 42'b100000001000010010000000000000000010001110;
    n1464[2003] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2002] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2001] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[2000] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1999] = 42'b100000000000000000000010000000000000000000;
    n1464[1998] = 42'b100000000000000000000010010000000000000000;
    n1464[1997] = 42'b000000000000000000000000000000000000000000;
    n1464[1996] = 42'b100000100000000000000000000000011010001100;
    n1464[1995] = 42'b000000000000000000000000000000000000000000;
    n1464[1994] = 42'b101000000000000000000000000000000000001110;
    n1464[1993] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1992] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1991] = 42'b100000000000000000000010000000000000000000;
    n1464[1990] = 42'b100000000000000000000010010000000000000000;
    n1464[1989] = 42'b000000000000000000000000000000000000000000;
    n1464[1988] = 42'b100000110111000000000000000000010000001100;
    n1464[1987] = 42'b000000000000000000000000000000000000000000;
    n1464[1986] = 42'b000000000000000000000000000000000000000000;
    n1464[1985] = 42'b101000000000000000000000000000000000001110;
    n1464[1984] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1983] = 42'b100000000000000000000010000000000000000000;
    n1464[1982] = 42'b100000000000000000000000000000000000000000;
    n1464[1981] = 42'b101010000000000000110000000000000000001010;
    n1464[1980] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1979] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1978] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1977] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1976] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1975] = 42'b100000000000000000000010000000000000000000;
    n1464[1974] = 42'b100000001000010010000010000000000010000010;
    n1464[1973] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1972] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1971] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1970] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1969] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1968] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1967] = 42'b100000000000000000000010000000000000000000;
    n1464[1966] = 42'b100000100000010010000000000000001010000010;
    n1464[1965] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1964] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1963] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1962] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1961] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1960] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1959] = 42'b100000000000000000000010000000000000000000;
    n1464[1958] = 42'b000000000000000000000000000000000000000010;
    n1464[1957] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1956] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1955] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1954] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1953] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1952] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1951] = 42'b100000000000000000000010000000000000000000;
    n1464[1950] = 42'b100000000000000000000010010000000000000000;
    n1464[1949] = 42'b100000000000000000000010000010000000000000;
    n1464[1948] = 42'b000000000000000000000000000000000000000000;
    n1464[1947] = 42'b100000111000010000000000000000011010000100;
    n1464[1946] = 42'b000000000000000000000000000000000000000000;
    n1464[1945] = 42'b101000000000000000000000000000000000000110;
    n1464[1944] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1943] = 42'b100000000000000000000010000000000000000000;
    n1464[1942] = 42'b100000000000000000000010010000000000000000;
    n1464[1941] = 42'b100000000000000000000010000010000000000000;
    n1464[1940] = 42'b000000000000000000000000000000000000000000;
    n1464[1939] = 42'b100000001000010010000000000000000010000110;
    n1464[1938] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1937] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1936] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1935] = 42'b100000000000000000000010000000000000000000;
    n1464[1934] = 42'b100000000000000000000010010000000000000000;
    n1464[1933] = 42'b100000000000000000000010000010000000000000;
    n1464[1932] = 42'b000000000000000000000000000000000000000000;
    n1464[1931] = 42'b100000100000000000000000000000011010000100;
    n1464[1930] = 42'b000000000000000000000000000000000000000000;
    n1464[1929] = 42'b101000000000000000000000000000000000000110;
    n1464[1928] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1927] = 42'b100000000000000000000010000000000000000000;
    n1464[1926] = 42'b100000000000000000000010010000000000000000;
    n1464[1925] = 42'b000000000000000000000000000000000000000000;
    n1464[1924] = 42'b000000000000000000000000000000000000000000;
    n1464[1923] = 42'b100000000000000000000000000000000000001100;
    n1464[1922] = 42'b100000000000000000000010010000000000000010;
    n1464[1921] = 42'b000000000000000000001000000000000000000000;
    n1464[1920] = 42'b000000000000000000000000000000000000000010;
    n1464[1919] = 42'b100000000000000000000010000000000000000000;
    n1464[1918] = 42'b100000000000000000000010010000000000000010;
    n1464[1917] = 42'b100000000000000000000000000000000000000000;
    n1464[1916] = 42'b000000000000000000001000000000000000000010;
    n1464[1915] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1914] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1913] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1912] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1911] = 42'b100000000000000000000010000000000000000000;
    n1464[1910] = 42'b100000000000000000000010010000000000000000;
    n1464[1909] = 42'b000000000000000000000000000000000000000000;
    n1464[1908] = 42'b100000000000000000000000100000000000001100;
    n1464[1907] = 42'b100000000000000000000001100010000000001100;
    n1464[1906] = 42'b100000000000000000000000000110000000000000;
    n1464[1905] = 42'b100000001000010010000000000000000010000110;
    n1464[1904] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1903] = 42'b100000000000000000000010000000000000000000;
    n1464[1902] = 42'b100000000000000000000010010000000000000000;
    n1464[1901] = 42'b000000000000000000000000000000000000000000;
    n1464[1900] = 42'b100000000000000000000000100000000000001100;
    n1464[1899] = 42'b100000000000000000000001010010000000001100;
    n1464[1898] = 42'b000000000000000000000000000000000000000000;
    n1464[1897] = 42'b100000001000010010000000000000000010000110;
    n1464[1896] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1895] = 42'b100000000000000000000010000000000000000000;
    n1464[1894] = 42'b100000000000000000000010000000010000000000;
    n1464[1893] = 42'b000000000000000000000000000000000000000000;
    n1464[1892] = 42'b101000000000000000000000000000000000010110;
    n1464[1891] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1890] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1889] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1888] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1887] = 42'b100000000000000000000010000000000000000000;
    n1464[1886] = 42'b100000000000000000000010010000000000000000;
    n1464[1885] = 42'b000000000000000000000000000000000000000000;
    n1464[1884] = 42'b100000110100010000000000000000011010001100;
    n1464[1883] = 42'b000000000000000000000000000000000000000000;
    n1464[1882] = 42'b101000000000000000000000000000000000001110;
    n1464[1881] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1880] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1879] = 42'b100000000000000000000010000000000000000000;
    n1464[1878] = 42'b100000000000000000000010010000000000000000;
    n1464[1877] = 42'b000000000000000000000000110000000000000000;
    n1464[1876] = 42'b100000001000010010000000000000000010001110;
    n1464[1875] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1874] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1873] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1872] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1871] = 42'b100000000000000000000010000000000000000000;
    n1464[1870] = 42'b100000000000000000000010010000000000000000;
    n1464[1869] = 42'b000000000000000000000000110000000000000000;
    n1464[1868] = 42'b100000100000000000000000000000011010001100;
    n1464[1867] = 42'b000000000000000000000000000000000000000000;
    n1464[1866] = 42'b101000000000000000000000000000000000001110;
    n1464[1865] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1864] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1863] = 42'b100000000000000000000010000000000000000000;
    n1464[1862] = 42'b100000000000000000000010010000000000000000;
    n1464[1861] = 42'b000000000000000000000000000000000000000000;
    n1464[1860] = 42'b100000110111000000000000000000010000001100;
    n1464[1859] = 42'b000000000000000000000000000000000000000000;
    n1464[1858] = 42'b000000000000000000000000000000000000000000;
    n1464[1857] = 42'b101000000000000000000000000000000000001110;
    n1464[1856] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1855] = 42'b100000000000000000000010000000000000000000;
    n1464[1854] = 42'b100000000000000000000000000000001000000010;
    n1464[1853] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1852] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1851] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1850] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1849] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1848] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1847] = 42'b100000000000000000000010000000000000000000;
    n1464[1846] = 42'b100000000000000000000010010000000000000000;
    n1464[1845] = 42'b100000000000000000000011000010000000000000;
    n1464[1844] = 42'b000000000000000000000000000110000000000000;
    n1464[1843] = 42'b100000001000010010000000000000000010000110;
    n1464[1842] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1841] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1840] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1839] = 42'b100000000000000000000010000000000000000000;
    n1464[1838] = 42'b100000011100010010000000000000000010000010;
    n1464[1837] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1836] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1835] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1834] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1833] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1832] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1831] = 42'b100000000000000000000010000000000000000000;
    n1464[1830] = 42'b000000000000000000000000000000000000000010;
    n1464[1829] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1828] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1827] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1826] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1825] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1824] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1823] = 42'b100000000000000000000010000000000000000000;
    n1464[1822] = 42'b100000000000000000000010010000000000000000;
    n1464[1821] = 42'b100000000000000000000010000010000000000000;
    n1464[1820] = 42'b000000000000000000000000000000000000000000;
    n1464[1819] = 42'b100000110100010000000000000000011010000100;
    n1464[1818] = 42'b000000000000000000000000000000000000000000;
    n1464[1817] = 42'b101000000000000000000000000000000000000110;
    n1464[1816] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1815] = 42'b100000000000000000000010000000000000000000;
    n1464[1814] = 42'b100000000000000000000010010000000000000000;
    n1464[1813] = 42'b100000000000000000000010110010000000000000;
    n1464[1812] = 42'b000000000000000000000000000110000000000000;
    n1464[1811] = 42'b100000001000010010000000000000000010000110;
    n1464[1810] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1809] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1808] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1807] = 42'b100000000000000000000010000000000000000000;
    n1464[1806] = 42'b100000000000000000000010010000000000000000;
    n1464[1805] = 42'b100000000000000000000010110010000000000000;
    n1464[1804] = 42'b000000000000000000000000000110000000000000;
    n1464[1803] = 42'b100000100000000000000000000000011010000100;
    n1464[1802] = 42'b000000000000000000000000000000000000000000;
    n1464[1801] = 42'b101000000000000000000000000000000000000110;
    n1464[1800] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1799] = 42'b100000000000000000000010000000000000000000;
    n1464[1798] = 42'b100000000000000000000010010000000000000000;
    n1464[1797] = 42'b000000000000000000000000000000000000000000;
    n1464[1796] = 42'b000000000000000000000000000000000000000000;
    n1464[1795] = 42'b100000000000000000000000000000000000001100;
    n1464[1794] = 42'b100000000000000000000010010000000000000010;
    n1464[1793] = 42'b000000000000000000001000000000000000000000;
    n1464[1792] = 42'b000000000000000000000000000000000000000010;
    n1464[1791] = 42'b100000000000000000000010000000000000000000;
    n1464[1790] = 42'b100000000000000000000010010000000000000000;
    n1464[1789] = 42'b100000000000000000000000000010000000000000;
    n1464[1788] = 42'b000000000000000000000000000000000000000000;
    n1464[1787] = 42'b101100000000000000110000000000000000001000;
    n1464[1786] = 42'b101110000000000000110000000000000000001000;
    n1464[1785] = 42'b000000000000000000001100000000000000000010;
    n1464[1784] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1783] = 42'b100000000000000000000010000000000000000000;
    n1464[1782] = 42'b100000000000000000000010010000000000000000;
    n1464[1781] = 42'b000000000000000000000000110000000000000000;
    n1464[1780] = 42'b100000000000000000000000100000000000001100;
    n1464[1779] = 42'b100000000000000000000001010010000000001100;
    n1464[1778] = 42'b000000000000000000000000000000000000000000;
    n1464[1777] = 42'b100000000100010010000000000000000010000110;
    n1464[1776] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1775] = 42'b100000000000000000000010000000000000000000;
    n1464[1774] = 42'b100000000000010100000000000000100000000000;
    n1464[1773] = 42'b000000000001010010000000000000000000000010;
    n1464[1772] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1771] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1770] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1769] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1768] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1767] = 42'b100000000000000000000010000000000000000000;
    n1464[1766] = 42'b100000000000000000000010000000010000000000;
    n1464[1765] = 42'b000000000000000000000000000000000000000000;
    n1464[1764] = 42'b101000000000000000000000000000000000010110;
    n1464[1763] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1762] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1761] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1760] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1759] = 42'b100000000000000000000010000000000000000000;
    n1464[1758] = 42'b100000000000000000000010010000000000000000;
    n1464[1757] = 42'b000000000000000000000000000000000000000000;
    n1464[1756] = 42'b100000110000010000000000000000001010001110;
    n1464[1755] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1754] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1753] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1752] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1751] = 42'b100000000000000000000010000000000000000000;
    n1464[1750] = 42'b100000000000000000000010010000000000000000;
    n1464[1749] = 42'b000000000000000000000000000000000000000000;
    n1464[1748] = 42'b100000000100010010000000000000000010001110;
    n1464[1747] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1746] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1745] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1744] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1743] = 42'b100000000000000000000010000000000000000000;
    n1464[1742] = 42'b100000000000000000000010010000000000000000;
    n1464[1741] = 42'b000000000000000000000000000000000000000000;
    n1464[1740] = 42'b100000101000000000000000000000011010001100;
    n1464[1739] = 42'b000000000000000000000000000000000000000000;
    n1464[1738] = 42'b101000000000000000000000000000000000001110;
    n1464[1737] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1736] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1735] = 42'b100000000000000000000010000000000000000000;
    n1464[1734] = 42'b100000000000000000000010010000000000000000;
    n1464[1733] = 42'b000000000000000000000000000000000000000000;
    n1464[1732] = 42'b100000110111000000000000000000010000001100;
    n1464[1731] = 42'b000000000000000000000000000000000000000000;
    n1464[1730] = 42'b000000000000000000000000000000000000000000;
    n1464[1729] = 42'b101000000000000000000000000000000000001110;
    n1464[1728] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1727] = 42'b100000000000000000000010000000000000000000;
    n1464[1726] = 42'b000000000000000000000000000000000000000000;
    n1464[1725] = 42'b000000000000000000100000000000000000000000;
    n1464[1724] = 42'b100000000000000000000000000000000110001010;
    n1464[1723] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1722] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1721] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1720] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1719] = 42'b100000000000000000000010000000000000000000;
    n1464[1718] = 42'b100000000100010010000010000000000010000010;
    n1464[1717] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1716] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1715] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1714] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1713] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1712] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1711] = 42'b100000000000000000000010000000000000000000;
    n1464[1710] = 42'b100000101000010010000000000000001010000010;
    n1464[1709] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1708] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1707] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1706] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1705] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1704] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1703] = 42'b100000000000000000000010000000000000000000;
    n1464[1702] = 42'b000000000000000000000000000000000000000010;
    n1464[1701] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1700] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1699] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1698] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1697] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1696] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1695] = 42'b100000000000000000000010000000000000000000;
    n1464[1694] = 42'b100000000000000000000010010000000000000000;
    n1464[1693] = 42'b100000000000000000000010000010000000000000;
    n1464[1692] = 42'b000000000000000000000000000000000000000000;
    n1464[1691] = 42'b100000110000010000000000000000001010000110;
    n1464[1690] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1689] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1688] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1687] = 42'b100000000000000000000010000000000000000000;
    n1464[1686] = 42'b100000000000000000000010010000000000000000;
    n1464[1685] = 42'b100000000000000000000010000010000000000000;
    n1464[1684] = 42'b000000000000000000000000000000000000000000;
    n1464[1683] = 42'b100000000100010010000000000000000010000110;
    n1464[1682] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1681] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1680] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1679] = 42'b100000000000000000000010000000000000000000;
    n1464[1678] = 42'b100000000000000000000010010000000000000000;
    n1464[1677] = 42'b100000000000000000000010000010000000000000;
    n1464[1676] = 42'b000000000000000000000000000000000000000000;
    n1464[1675] = 42'b100000101000000000000000000000011010000100;
    n1464[1674] = 42'b000000000000000000000000000000000000000000;
    n1464[1673] = 42'b101000000000000000000000000000000000000110;
    n1464[1672] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1671] = 42'b100000000000000000000010000000000000000000;
    n1464[1670] = 42'b100000000000000000000010010000000000000000;
    n1464[1669] = 42'b000000000000000000000000000000000000000000;
    n1464[1668] = 42'b000000000000000000000000000000000000000000;
    n1464[1667] = 42'b100000000000000000000000000000000000001100;
    n1464[1666] = 42'b100000000000000000000010010000000000000010;
    n1464[1665] = 42'b000000000000000000001000000000000000000000;
    n1464[1664] = 42'b000000000000000000000000000000000000000010;
    n1464[1663] = 42'b100000000000000000000010000000000000000000;
    n1464[1662] = 42'b100000000000000000000010010000000000000010;
    n1464[1661] = 42'b100000000000000000000000000000000000000000;
    n1464[1660] = 42'b000000000000000000001000000000000000000010;
    n1464[1659] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1658] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1657] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1656] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1655] = 42'b100000000000000000000010000000000000000000;
    n1464[1654] = 42'b100000000000000000000010010000000000000000;
    n1464[1653] = 42'b000000000000000000000000000000000000000000;
    n1464[1652] = 42'b100000000000000000000000100000000000001100;
    n1464[1651] = 42'b100000000000000000000001100010000000001100;
    n1464[1650] = 42'b000000000000000000000000000110000000000000;
    n1464[1649] = 42'b100000000100010010000000000000000010000110;
    n1464[1648] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1647] = 42'b100000000000000000000010000000000000000000;
    n1464[1646] = 42'b100000000000000000000010010000000000000000;
    n1464[1645] = 42'b000000000000000000000000000000000000000000;
    n1464[1644] = 42'b100000000000000000000000100000000000001100;
    n1464[1643] = 42'b100000000000000000000001010010000000001100;
    n1464[1642] = 42'b000000000000000000000000000000000000000000;
    n1464[1641] = 42'b100000000100010010000000000000000010000110;
    n1464[1640] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1639] = 42'b100000000000000000000010000000000000000000;
    n1464[1638] = 42'b000000000000000000000000000000000000000010;
    n1464[1637] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1636] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1635] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1634] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1633] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1632] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1631] = 42'b100000000000000000000010000000000000000000;
    n1464[1630] = 42'b100000000000000000000010010000000000000000;
    n1464[1629] = 42'b000000000000000000000000110000000000000000;
    n1464[1628] = 42'b100000110000010000000000000000001010001110;
    n1464[1627] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1626] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1625] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1624] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1623] = 42'b100000000000000000000010000000000000000000;
    n1464[1622] = 42'b100000000000000000000010010000000000000000;
    n1464[1621] = 42'b000000000000000000000000110000000000000000;
    n1464[1620] = 42'b100000000100010010000000000000000010001110;
    n1464[1619] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1618] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1617] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1616] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1615] = 42'b100000000000000000000010000000000000000000;
    n1464[1614] = 42'b100000000000000000000010010000000000000000;
    n1464[1613] = 42'b000000000000000000000000110000000000000000;
    n1464[1612] = 42'b100000101000000000000000000000011010001100;
    n1464[1611] = 42'b000000000000000000000000000000000000000000;
    n1464[1610] = 42'b101000000000000000000000000000000000001110;
    n1464[1609] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1608] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1607] = 42'b100000000000000000000010000000000000000000;
    n1464[1606] = 42'b100000000000000000000010010000000000000000;
    n1464[1605] = 42'b000000000000000000000000000000000000000000;
    n1464[1604] = 42'b100000110111000000000000000000010000001100;
    n1464[1603] = 42'b000000000000000000000000000000000000000000;
    n1464[1602] = 42'b000000000000000000000000000000000000000000;
    n1464[1601] = 42'b101000000000000000000000000000000000001110;
    n1464[1600] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1599] = 42'b100000000000000000000010000000000000000000;
    n1464[1598] = 42'b100000000000000000000000000000001000000010;
    n1464[1597] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1596] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1595] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1594] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1593] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1592] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1591] = 42'b100000000000000000000010000000000000000000;
    n1464[1590] = 42'b100000000000000000000010010000000000000000;
    n1464[1589] = 42'b100000000000000000000011000010000000000000;
    n1464[1588] = 42'b000000000000000000000000000110000000000000;
    n1464[1587] = 42'b100000000100010010000000000000000010000110;
    n1464[1586] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1585] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1584] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1583] = 42'b100000000000000000000010000000000000000000;
    n1464[1582] = 42'b100000011000010010000000000000000010000010;
    n1464[1581] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1580] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1579] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1578] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1577] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1576] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1575] = 42'b100000000000000000000010000000000000000000;
    n1464[1574] = 42'b000000000000000000000000000000000000000010;
    n1464[1573] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1572] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1571] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1570] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1569] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1568] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1567] = 42'b100000000000000000000010000000000000000000;
    n1464[1566] = 42'b100000000000000000000010010000000000000000;
    n1464[1565] = 42'b100000000000000000000010110010000000000000;
    n1464[1564] = 42'b000000000000000000000000000110000000000000;
    n1464[1563] = 42'b100000110000010000000000000000001010000110;
    n1464[1562] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1561] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1560] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1559] = 42'b100000000000000000000010000000000000000000;
    n1464[1558] = 42'b100000000000000000000010010000000000000000;
    n1464[1557] = 42'b100000000000000000000010110010000000000000;
    n1464[1556] = 42'b000000000000000000000000000110000000000000;
    n1464[1555] = 42'b100000000100010010000000000000000010000110;
    n1464[1554] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1553] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1552] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1551] = 42'b100000000000000000000010000000000000000000;
    n1464[1550] = 42'b100000000000000000000010010000000000000000;
    n1464[1549] = 42'b100000000000000000000010110010000000000000;
    n1464[1548] = 42'b000000000000000000000000000110000000000000;
    n1464[1547] = 42'b100000101000000000000000000000011010000100;
    n1464[1546] = 42'b000000000000000000000000000000000000000000;
    n1464[1545] = 42'b101000000000000000000000000000000000000110;
    n1464[1544] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1543] = 42'b100000000000000000000010000000000000000000;
    n1464[1542] = 42'b100000000000000000000010010000000000000000;
    n1464[1541] = 42'b000000000000000000000000000000000000000000;
    n1464[1540] = 42'b000000000000000000000000000000000000000000;
    n1464[1539] = 42'b100000000000000000000000000000000000001100;
    n1464[1538] = 42'b100000000000000000000010010000000000000010;
    n1464[1537] = 42'b000000000000000000001000000000000000000000;
    n1464[1536] = 42'b000000000000000000000000000000000000000010;
    n1464[1535] = 42'b100000000000000000000010000000000000000000;
    n1464[1534] = 42'b000000000000000000000000000000000000000000;
    n1464[1533] = 42'b000000000000000000000000000000000000000000;
    n1464[1532] = 42'b000000000000000000100000000000000000000000;
    n1464[1531] = 42'b100000000000000000100000000000000110001000;
    n1464[1530] = 42'b100000000000000000100100000000000000001000;
    n1464[1529] = 42'b100000000000000000000110000000000000001010;
    n1464[1528] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1527] = 42'b100000000000000000000010000000000000000000;
    n1464[1526] = 42'b100000000000000000000010010000000000000000;
    n1464[1525] = 42'b000000000000000000000000110000000000000000;
    n1464[1524] = 42'b100000000000000000000000100000000000001100;
    n1464[1523] = 42'b100000000000000000000001010010000000001100;
    n1464[1522] = 42'b000000000000000000000000000000000000000000;
    n1464[1521] = 42'b100000001100010010000000000000000010000110;
    n1464[1520] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1519] = 42'b100000000000000000000010000000000000000000;
    n1464[1518] = 42'b100000000001001000000000000000110000000000;
    n1464[1517] = 42'b000000000001000010000000000000000000000010;
    n1464[1516] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1515] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1514] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1513] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1512] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1511] = 42'b100000000000000000000010000000000000000000;
    n1464[1510] = 42'b100000000000000000000010000000010000000000;
    n1464[1509] = 42'b000000000000000000000000000000000000000000;
    n1464[1508] = 42'b000000000010110010000000000000000000000010;
    n1464[1507] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1506] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1505] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1504] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1503] = 42'b100000000000000000000010000000000000000000;
    n1464[1502] = 42'b000000000000000000000000000000000000000000;
    n1464[1501] = 42'b101100000000000000110000000000000000001000;
    n1464[1500] = 42'b101110000000000000110000000000000000001000;
    n1464[1499] = 42'b100000000000000000000010010000000000000000;
    n1464[1498] = 42'b000000000000000000000000000000000000000000;
    n1464[1497] = 42'b000000000000000000000000000000000000000000;
    n1464[1496] = 42'b000000000000000000001000000000000000000010;
    n1464[1495] = 42'b100000000000000000000010000000000000000000;
    n1464[1494] = 42'b100000000000000000000010010000000000000000;
    n1464[1493] = 42'b000000000000000000000000000000000000000000;
    n1464[1492] = 42'b100000001100010010000000000000000010001110;
    n1464[1491] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1490] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1489] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1488] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1487] = 42'b100000000000000000000010000000000000000000;
    n1464[1486] = 42'b100000000000000000000010010000000000000000;
    n1464[1485] = 42'b000000000000000000000000000000000000000000;
    n1464[1484] = 42'b100000100100000000000000000000011010001100;
    n1464[1483] = 42'b000000000000000000000000000000000000000000;
    n1464[1482] = 42'b101000000000000000000000000000000000001110;
    n1464[1481] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1480] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1479] = 42'b100000000000000000000010000000000000000000;
    n1464[1478] = 42'b100000000000000000000010010000000000000000;
    n1464[1477] = 42'b000000000000000000000000000000000000000000;
    n1464[1476] = 42'b100000110111000000000000000000010000001100;
    n1464[1475] = 42'b000000000000000000000000000000000000000000;
    n1464[1474] = 42'b000000000000000000000000000000000000000000;
    n1464[1473] = 42'b101000000000000000000000000000000000001110;
    n1464[1472] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1471] = 42'b100000000000000000000010000000000000000000;
    n1464[1470] = 42'b100000000000000000000000000000000000000000;
    n1464[1469] = 42'b100010000000000000110000000000000000001010;
    n1464[1468] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1467] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1466] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1465] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1464] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1463] = 42'b100000000000000000000010000000000000000000;
    n1464[1462] = 42'b100000001100010010000010000000000010000010;
    n1464[1461] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1460] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1459] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1458] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1457] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1456] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1455] = 42'b100000000000000000000010000000000000000000;
    n1464[1454] = 42'b100000100100010010000000000000001010000010;
    n1464[1453] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1452] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1451] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1450] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1449] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1448] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1447] = 42'b100000000000000000000010000000000000000000;
    n1464[1446] = 42'b000000000000000000000000000000000000000010;
    n1464[1445] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1444] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1443] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1442] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1441] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1440] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1439] = 42'b100000000000000000000010000000000000000000;
    n1464[1438] = 42'b100000000000000000000010010000000000000000;
    n1464[1437] = 42'b100000000000000000000000000010000000000000;
    n1464[1436] = 42'b000000000000000000001100000000000000000010;
    n1464[1435] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1434] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1433] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1432] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1431] = 42'b100000000000000000000010000000000000000000;
    n1464[1430] = 42'b100000000000000000000010010000000000000000;
    n1464[1429] = 42'b100000000000000000000010000010000000000000;
    n1464[1428] = 42'b000000000000000000000000000000000000000000;
    n1464[1427] = 42'b100000001100010010000000000000000010000110;
    n1464[1426] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1425] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1424] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1423] = 42'b100000000000000000000010000000000000000000;
    n1464[1422] = 42'b100000000000000000000010010000000000000000;
    n1464[1421] = 42'b100000000000000000000010000010000000000000;
    n1464[1420] = 42'b000000000000000000000000000000000000000000;
    n1464[1419] = 42'b100000100100000000000000000000011010000100;
    n1464[1418] = 42'b000000000000000000000000000000000000000000;
    n1464[1417] = 42'b101000000000000000000000000000000000000110;
    n1464[1416] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1415] = 42'b100000000000000000000010000000000000000000;
    n1464[1414] = 42'b100000000000000000000010010000000000000000;
    n1464[1413] = 42'b000000000000000000000000000000000000000000;
    n1464[1412] = 42'b000000000000000000000000000000000000000000;
    n1464[1411] = 42'b100000000000000000000000000000000000001100;
    n1464[1410] = 42'b100000000000000000000010010000000000000010;
    n1464[1409] = 42'b000000000000000000001000000000000000000000;
    n1464[1408] = 42'b000000000000000000000000000000000000000010;
    n1464[1407] = 42'b100000000000000000000010000000000000000000;
    n1464[1406] = 42'b100000000000000000000010010000000000000010;
    n1464[1405] = 42'b100000000000000000000000000000000000000000;
    n1464[1404] = 42'b000000000000000000001000000000000000000010;
    n1464[1403] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1402] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1401] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1400] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1399] = 42'b100000000000000000000010000000000000000000;
    n1464[1398] = 42'b100000000000000000000010010000000000000000;
    n1464[1397] = 42'b000000000000000000000000000000000000000000;
    n1464[1396] = 42'b100000000000000000000000100000000000001100;
    n1464[1395] = 42'b100000000000000000000001100010000000001100;
    n1464[1394] = 42'b000000000000000000000000000110000000000000;
    n1464[1393] = 42'b100000001100010010000000000000000010000110;
    n1464[1392] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1391] = 42'b100000000000000000000010000000000000000000;
    n1464[1390] = 42'b100000000000000000000010010000000000000000;
    n1464[1389] = 42'b000000000000000000000000000000000000000000;
    n1464[1388] = 42'b100000000000000000000000100000000000001100;
    n1464[1387] = 42'b100000000000000000000001010010000000001100;
    n1464[1386] = 42'b000000000000000000000000000000000000000000;
    n1464[1385] = 42'b100000001100010010000000000000000010000110;
    n1464[1384] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1383] = 42'b100000000000000000000010000000000000000000;
    n1464[1382] = 42'b100000000000000000000010000000010000000000;
    n1464[1381] = 42'b000000000000000000000000000000000000000000;
    n1464[1380] = 42'b000000000000000000000000000000000000000000;
    n1464[1379] = 42'b000000000000000000000000000000000000000010;
    n1464[1378] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1377] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1376] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1375] = 42'b100000000000000000000010000000000000000000;
    n1464[1374] = 42'b100000000000000000000000000000000000000000;
    n1464[1373] = 42'b000000000000000000000000000000000000000010;
    n1464[1372] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1371] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1370] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1369] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1368] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1367] = 42'b100000000000000000000010000000000000000000;
    n1464[1366] = 42'b100000000000000000000010010000000000000000;
    n1464[1365] = 42'b000000000000000000000000110000000000000000;
    n1464[1364] = 42'b100000001100010010000000000000000010001110;
    n1464[1363] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1362] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1361] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1360] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1359] = 42'b100000000000000000000010000000000000000000;
    n1464[1358] = 42'b100000000000000000000010010000000000000000;
    n1464[1357] = 42'b000000000000000000000000110000000000000000;
    n1464[1356] = 42'b100000100100000000000000000000011010001100;
    n1464[1355] = 42'b000000000000000000000000000000000000000000;
    n1464[1354] = 42'b101000000000000000000000000000000000001110;
    n1464[1353] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1352] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1351] = 42'b100000000000000000000010000000000000000000;
    n1464[1350] = 42'b100000000000000000000010010000000000000000;
    n1464[1349] = 42'b000000000000000000000000000000000000000000;
    n1464[1348] = 42'b100000110111000000000000000000010000001100;
    n1464[1347] = 42'b000000000000000000000000000000000000000000;
    n1464[1346] = 42'b000000000000000000000000000000000000000000;
    n1464[1345] = 42'b101000000000000000000000000000000000001110;
    n1464[1344] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1343] = 42'b100000000000000000000010000000000000000000;
    n1464[1342] = 42'b100000000000000000000000000000001000000010;
    n1464[1341] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1340] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1339] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1338] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1337] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1336] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1335] = 42'b100000000000000000000010000000000000000000;
    n1464[1334] = 42'b100000000000000000000010010000000000000000;
    n1464[1333] = 42'b100000000000000000000011000010000000000000;
    n1464[1332] = 42'b000000000000000000000000000110000000000000;
    n1464[1331] = 42'b100000001100010010000000000000000010000110;
    n1464[1330] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1329] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1328] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1327] = 42'b100000000000000000000010000000000000000000;
    n1464[1326] = 42'b100000000000000000000000000000000000000000;
    n1464[1325] = 42'b100110000000000000110000000000000000001010;
    n1464[1324] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1323] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1322] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1321] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1320] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1319] = 42'b100000000000000000000010000000000000000000;
    n1464[1318] = 42'b000000000000000000000000000000000000000010;
    n1464[1317] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1316] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1315] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1314] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1313] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1312] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1311] = 42'b100000000000000000000010000000000000000000;
    n1464[1310] = 42'b000000000000000000000000000000000000000010;
    n1464[1309] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1308] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1307] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1306] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1305] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1304] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1303] = 42'b100000000000000000000010000000000000000000;
    n1464[1302] = 42'b100000000000000000000010010000000000000000;
    n1464[1301] = 42'b100000000000000000000010110010000000000000;
    n1464[1300] = 42'b000000000000000000000000000110000000000000;
    n1464[1299] = 42'b100000001100010010000000000000000010000110;
    n1464[1298] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1297] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1296] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1295] = 42'b100000000000000000000010000000000000000000;
    n1464[1294] = 42'b100000000000000000000010010000000000000000;
    n1464[1293] = 42'b100000000000000000000010110010000000000000;
    n1464[1292] = 42'b000000000000000000000000000110000000000000;
    n1464[1291] = 42'b100000100100000000000000000000011010000100;
    n1464[1290] = 42'b000000000000000000000000000000000000000000;
    n1464[1289] = 42'b101000000000000000000000000000000000000110;
    n1464[1288] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1287] = 42'b100000000000000000000010000000000000000000;
    n1464[1286] = 42'b100000000000000000000010010000000000000000;
    n1464[1285] = 42'b000000000000000000000000000000000000000000;
    n1464[1284] = 42'b000000000000000000000000000000000000000000;
    n1464[1283] = 42'b100000000000000000000000000000000000001100;
    n1464[1282] = 42'b100000000000000000000010010000000000000010;
    n1464[1281] = 42'b000000000000000000001000000000000000000000;
    n1464[1280] = 42'b000000000000000000000000000000000000000010;
    n1464[1279] = 42'b100000000000000000000010000000000000000000;
    n1464[1278] = 42'b000000000000000000000000000000000000000000;
    n1464[1277] = 42'b000000000000000000000000000000000000000000;
    n1464[1276] = 42'b000000000000000000100000000000000000000000;
    n1464[1275] = 42'b100000000000000000100100000000000000001000;
    n1464[1274] = 42'b100000000000000000000110000000000000001000;
    n1464[1273] = 42'b000000000000000000000010000000000000000010;
    n1464[1272] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1271] = 42'b100000000000000000000010000000000000000000;
    n1464[1270] = 42'b100000000000000000000010010000000000000000;
    n1464[1269] = 42'b000000000000000000000000110000000000000000;
    n1464[1268] = 42'b100000000000000000000000100000000000001100;
    n1464[1267] = 42'b100000000000000000000001010010000000001100;
    n1464[1266] = 42'b000000000000000000000000000000000000000000;
    n1464[1265] = 42'b100000010000010010000000000000001010000101;
    n1464[1264] = 42'b100000000000000000000000000000000000000010;
    n1464[1263] = 42'b100000000000000000000010000000000000000000;
    n1464[1262] = 42'b100000000011110010000000000000000000000010;
    n1464[1261] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1260] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1259] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1258] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1257] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1256] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1255] = 42'b100000000000000000000010000000000000000000;
    n1464[1254] = 42'b000000000000000000000000000000000000000010;
    n1464[1253] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1252] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1251] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1250] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1249] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1248] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1247] = 42'b100000000000000000000010000000000000000000;
    n1464[1246] = 42'b100000000000000000000010010000000000000000;
    n1464[1245] = 42'b000000000000000000000000000000000000000000;
    n1464[1244] = 42'b111110000000000000000000000000000000001110;
    n1464[1243] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1242] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1241] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1240] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1239] = 42'b100000000000000000000010000000000000000000;
    n1464[1238] = 42'b100000000000000000000010010000000000000000;
    n1464[1237] = 42'b000000000000000000000000000000000000000000;
    n1464[1236] = 42'b100000010000010010000000000000001010001101;
    n1464[1235] = 42'b000000000000000000000000000000000000000010;
    n1464[1234] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1233] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1232] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1231] = 42'b100000000000000000000010000000000000000000;
    n1464[1230] = 42'b100000000000000000000010010000000000000000;
    n1464[1229] = 42'b000000000000000000000000000000000000000000;
    n1464[1228] = 42'b100000101100000000000000000000011010001100;
    n1464[1227] = 42'b000000000000000000000000000000000000000000;
    n1464[1226] = 42'b101000000000000000000000000000000000001110;
    n1464[1225] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1224] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1223] = 42'b100000000000000000000010000000000000000000;
    n1464[1222] = 42'b100000000000000000000010010000000000000000;
    n1464[1221] = 42'b000000000000000000000000000000000000000000;
    n1464[1220] = 42'b100000110111000000000000000000010000001100;
    n1464[1219] = 42'b000000000000000000000000000000000000000000;
    n1464[1218] = 42'b000000000000000000000000000000000000000000;
    n1464[1217] = 42'b101000000000000000000000000000000000001110;
    n1464[1216] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1215] = 42'b100000000000000000000010000000000000000000;
    n1464[1214] = 42'b000000000000000000000000000000000000000000;
    n1464[1213] = 42'b000000000000000000100000000000000000000000;
    n1464[1212] = 42'b100000000000000010000000000000000010001010;
    n1464[1211] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1210] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1209] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1208] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1207] = 42'b100000000000000000000010000000000000000000;
    n1464[1206] = 42'b100000010000010010000010000000001010000001;
    n1464[1205] = 42'b000000000000000000000000000000000000000010;
    n1464[1204] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1203] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1202] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1201] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1200] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1199] = 42'b100000000000000000000010000000000000000000;
    n1464[1198] = 42'b100000101100010010000000000000001010000010;
    n1464[1197] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1196] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1195] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1194] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1193] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1192] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1191] = 42'b100000000000000000000010000000000000000000;
    n1464[1190] = 42'b000000000000000000000000000000000000000010;
    n1464[1189] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1188] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1187] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1186] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1185] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1184] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1183] = 42'b100000000000000000000010000000000000000000;
    n1464[1182] = 42'b100000000000000000000010010000000000000000;
    n1464[1181] = 42'b100000000000000000000010000010000000000000;
    n1464[1180] = 42'b000000000000000000000000000000000000000000;
    n1464[1179] = 42'b100000000000000000000100100000000000000100;
    n1464[1178] = 42'b000000000000000000000000000110000000000000;
    n1464[1177] = 42'b100000000000000000000110000000000000000110;
    n1464[1176] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1175] = 42'b100000000000000000000010000000000000000000;
    n1464[1174] = 42'b100000000000000000000010010000000000000000;
    n1464[1173] = 42'b100000000000000000000010000010000000000000;
    n1464[1172] = 42'b000000000000000000000000000000000000000000;
    n1464[1171] = 42'b100000010000010010000000000000001010000101;
    n1464[1170] = 42'b000000000000000000000000000000000000000010;
    n1464[1169] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1168] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1167] = 42'b100000000000000000000010000000000000000000;
    n1464[1166] = 42'b100000000000000000000010010000000000000000;
    n1464[1165] = 42'b100000000000000000000010000010000000000000;
    n1464[1164] = 42'b000000000000000000000000000000000000000000;
    n1464[1163] = 42'b100000101100000000000000000000011010000100;
    n1464[1162] = 42'b000000000000000000000000000000000000000000;
    n1464[1161] = 42'b101000000000000000000000000000000000000110;
    n1464[1160] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1159] = 42'b100000000000000000000010000000000000000000;
    n1464[1158] = 42'b100000000000000000000010010000000000000000;
    n1464[1157] = 42'b000000000000000000000000000000000000000000;
    n1464[1156] = 42'b000000000000000000000000000000000000000000;
    n1464[1155] = 42'b100000000000000000000000000000000000001100;
    n1464[1154] = 42'b100000000000000000000010010000000000000010;
    n1464[1153] = 42'b000000000000000000001000000000000000000000;
    n1464[1152] = 42'b000000000000000000000000000000000000000010;
    n1464[1151] = 42'b100000000000000000000010000000000000000000;
    n1464[1150] = 42'b100000000000000000000010010000000000000010;
    n1464[1149] = 42'b100000000000000000000000000000000000000000;
    n1464[1148] = 42'b000000000000000000001000000000000000000010;
    n1464[1147] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1146] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1145] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1144] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1143] = 42'b100000000000000000000010000000000000000000;
    n1464[1142] = 42'b100000000000000000000010010000000000000000;
    n1464[1141] = 42'b000000000000000000000000000000000000000000;
    n1464[1140] = 42'b100000000000000000000000100000000000001100;
    n1464[1139] = 42'b100000000000000000000001100010000000001100;
    n1464[1138] = 42'b000000000000000000000000000110000000000000;
    n1464[1137] = 42'b100000010000010010000000000000001010000101;
    n1464[1136] = 42'b000000000000000000000000000000000000000010;
    n1464[1135] = 42'b100000000000000000000010000000000000000000;
    n1464[1134] = 42'b100000000000000000000010010000000000000000;
    n1464[1133] = 42'b000000000000000000000000000000000000000000;
    n1464[1132] = 42'b100000000000000000000000100000000000001100;
    n1464[1131] = 42'b100000000000000000000001010010000000001100;
    n1464[1130] = 42'b000000000000000000000000000000000000000000;
    n1464[1129] = 42'b100000010000010010000000000000001010000101;
    n1464[1128] = 42'b000000000000000000000000000000000000000010;
    n1464[1127] = 42'b100000000000000000000010000000000000000000;
    n1464[1126] = 42'b100110000000000000110000000000000000001000;
    n1464[1125] = 42'b100010000000000000110000000000000000001000;
    n1464[1124] = 42'b100100000000000000000000000000000000001000;
    n1464[1123] = 42'b100000000000000100000010000000000000000000;
    n1464[1122] = 42'b100000000000000000000010000000000000100000;
    n1464[1121] = 42'b100000000000001000000010000000000000000000;
    n1464[1120] = 42'b100000000000000000000010000000000001000000;
    n1464[1119] = 42'b100000000000000000000010000000000000000000;
    n1464[1118] = 42'b100000000000000000000010010000000000000000;
    n1464[1117] = 42'b000000000000000000000000110000000000000000;
    n1464[1116] = 42'b111110000000000000000000000000000000001110;
    n1464[1115] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1114] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1113] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1112] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1111] = 42'b100000000000000000000010000000000000000000;
    n1464[1110] = 42'b100000000000000000000010010000000000000000;
    n1464[1109] = 42'b000000000000000000000000110000000000000000;
    n1464[1108] = 42'b100000010000010010000000000000001010001101;
    n1464[1107] = 42'b000000000000000000000000000000000000000010;
    n1464[1106] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1105] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1104] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1103] = 42'b100000000000000000000010000000000000000000;
    n1464[1102] = 42'b100000000000000000000010010000000000000000;
    n1464[1101] = 42'b000000000000000000000000110000000000000000;
    n1464[1100] = 42'b100000101100000000000000000000011010001100;
    n1464[1099] = 42'b000000000000000000000000000000000000000000;
    n1464[1098] = 42'b101000000000000000000000000000000000001110;
    n1464[1097] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1096] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1095] = 42'b100000000000000000000010000000000000000000;
    n1464[1094] = 42'b100000000000000000000010010000000000000000;
    n1464[1093] = 42'b000000000000000000000000000000000000000000;
    n1464[1092] = 42'b100000110111000000000000000000010000001100;
    n1464[1091] = 42'b000000000000000000000000000000000000000000;
    n1464[1090] = 42'b000000000000000000000000000000000000000000;
    n1464[1089] = 42'b101000000000000000000000000000000000001110;
    n1464[1088] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1087] = 42'b100000000000000000000010000000000000000000;
    n1464[1086] = 42'b100000000000000000000000000000001000000010;
    n1464[1085] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1084] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1083] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1082] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1081] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1080] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1079] = 42'b100000000000000000000010000000000000000000;
    n1464[1078] = 42'b100000000000000000000010010000000000000000;
    n1464[1077] = 42'b100000000000000000000011000010000000000000;
    n1464[1076] = 42'b000000000000000000000000000110000000000000;
    n1464[1075] = 42'b100000010000010010000000000000001010000101;
    n1464[1074] = 42'b000000000000000000000000000000000000000010;
    n1464[1073] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1072] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1071] = 42'b100000000000000000000010000000000000000000;
    n1464[1070] = 42'b000000000000000000000000000000000000000000;
    n1464[1069] = 42'b000000000000000000100000000000000000000000;
    n1464[1068] = 42'b100000000000001000000000000000000010001010;
    n1464[1067] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1066] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1065] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1064] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1063] = 42'b100000000000000000000010000000000000000000;
    n1464[1062] = 42'b000000000000000000000000000000000000000010;
    n1464[1061] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1060] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1059] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1058] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1057] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1056] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1055] = 42'b100000000000000000000010000000000000000000;
    n1464[1054] = 42'b100000000000000000000010010000000000000000;
    n1464[1053] = 42'b100000000000000000000010110010000000000000;
    n1464[1052] = 42'b000000000000000000000000000110000000000000;
    n1464[1051] = 42'b100000000000000000000100100000000000000100;
    n1464[1050] = 42'b000000000000000000000000000110000000000000;
    n1464[1049] = 42'b100000000000000000000110000000000000000110;
    n1464[1048] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1047] = 42'b100000000000000000000010000000000000000000;
    n1464[1046] = 42'b100000000000000000000010010000000000000000;
    n1464[1045] = 42'b100000000000000000000010110010000000000000;
    n1464[1044] = 42'b000000000000000000000000000110000000000000;
    n1464[1043] = 42'b100000010000010010000000000000001010000101;
    n1464[1042] = 42'b000000000000000000000000000000000000000010;
    n1464[1041] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1040] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1039] = 42'b100000000000000000000010000000000000000000;
    n1464[1038] = 42'b100000000000000000000010010000000000000000;
    n1464[1037] = 42'b100000000000000000000010110010000000000000;
    n1464[1036] = 42'b000000000000000000000000000110000000000000;
    n1464[1035] = 42'b100000101100000000000000000000011010000100;
    n1464[1034] = 42'b000000000000000000000000000000000000000000;
    n1464[1033] = 42'b101000000000000000000000000000000000000110;
    n1464[1032] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1031] = 42'b100000000000000000000010000000000000000000;
    n1464[1030] = 42'b100000000000000000000010010000000000000000;
    n1464[1029] = 42'b000000000000000000000000000000000000000000;
    n1464[1028] = 42'b000000000000000000000000000000000000000000;
    n1464[1027] = 42'b100000000000000000000000000000000000001100;
    n1464[1026] = 42'b100000000000000000000010010000000000000010;
    n1464[1025] = 42'b100000000000000000001000000000000000000000;
    n1464[1024] = 42'b000000000000000000000000000000000000000010;
    n1464[1023] = 42'b100000000000000000000010000000000000000000;
    n1464[1022] = 42'b100000000000000000000010010000000000000000;
    n1464[1021] = 42'b000000000000000000000000000000000000000000;
    n1464[1020] = 42'b000000000000000000001000000000000000000010;
    n1464[1019] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1018] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1017] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1016] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1015] = 42'b100000000000000000000010000000000000000000;
    n1464[1014] = 42'b100000000000000000000010010000000000000000;
    n1464[1013] = 42'b000000000000000000000000110000000000000000;
    n1464[1012] = 42'b100000000000000000000000100000000000001100;
    n1464[1011] = 42'b100000000000000000000001010010000000001100;
    n1464[1010] = 42'b000000000000000000000000000000000000000000;
    n1464[1009] = 42'b100010000000000000000000000000000000000110;
    n1464[1008] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1007] = 42'b100000000000000000000010000000000000000000;
    n1464[1006] = 42'b100000000011110100000000000000000000000010;
    n1464[1005] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1004] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1003] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1002] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1001] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[1000] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[999] = 42'b100000000000000000000010000000000000000000;
    n1464[998] = 42'b100000000000000000000010000000010000000000;
    n1464[997] = 42'b100000000000000000000010010000000000000000;
    n1464[996] = 42'b000000000000000000000000000000000000000000;
    n1464[995] = 42'b000000000000000000000000000000000000000000;
    n1464[994] = 42'b000000000000000000000000000000000000000000;
    n1464[993] = 42'b100000110001010000000000000000001010001110;
    n1464[992] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[991] = 42'b100000000000000000000010000000000000000000;
    n1464[990] = 42'b100000000000000000000010010000000000000000;
    n1464[989] = 42'b000000000000000000000000000000000000000000;
    n1464[988] = 42'b100110000000000000000000000000000000001110;
    n1464[987] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[986] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[985] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[984] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[983] = 42'b100000000000000000000010000000000000000000;
    n1464[982] = 42'b100000000000000000000010010000000000000000;
    n1464[981] = 42'b000000000000000000000000000000000000000000;
    n1464[980] = 42'b100010000000000000000000000000000000001110;
    n1464[979] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[978] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[977] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[976] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[975] = 42'b100000000000000000000010000000000000000000;
    n1464[974] = 42'b100000000000000000000010010000000000000000;
    n1464[973] = 42'b000000000000000000000000000000000000000000;
    n1464[972] = 42'b100100000000000000000000000000000000001110;
    n1464[971] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[970] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[969] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[968] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[967] = 42'b100000000000000000000010000000000000000000;
    n1464[966] = 42'b100000000000000000000010010000000000000000;
    n1464[965] = 42'b000000000000000000000000000000000000000000;
    n1464[964] = 42'b100000111011000000000000000000010000001100;
    n1464[963] = 42'b000000000000000000000000000000000000000000;
    n1464[962] = 42'b000000000000000000000000000000000000000000;
    n1464[961] = 42'b101000000000000000000000000000000000001110;
    n1464[960] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[959] = 42'b100000000000000000000010000000000000000000;
    n1464[958] = 42'b100000011000111000000000000000000010000010;
    n1464[957] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[956] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[955] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[954] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[953] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[952] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[951] = 42'b100000000000000000000010000000000000000000;
    n1464[950] = 42'b100000110000010000000010000000001010000010;
    n1464[949] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[948] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[947] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[946] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[945] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[944] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[943] = 42'b100000000000000000000010000000000000000000;
    n1464[942] = 42'b100000000000100010000000000000000010000010;
    n1464[941] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[940] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[939] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[938] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[937] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[936] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[935] = 42'b100000000000000000000010000000000000000000;
    n1464[934] = 42'b000000000000000000000000000000000000000010;
    n1464[933] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[932] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[931] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[930] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[929] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[928] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[927] = 42'b100000000000000000000010000000000000000000;
    n1464[926] = 42'b100000000000000000000010010000000000000000;
    n1464[925] = 42'b100000000000000000000010000010000000000000;
    n1464[924] = 42'b000000000000000000000000000000000000000000;
    n1464[923] = 42'b100110000000000000000000000000000000000110;
    n1464[922] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[921] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[920] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[919] = 42'b100000000000000000000010000000000000000000;
    n1464[918] = 42'b100000000000000000000010010000000000000000;
    n1464[917] = 42'b100000000000000000000010000010000000000000;
    n1464[916] = 42'b000000000000000000000000000000000000000000;
    n1464[915] = 42'b100010000000000000000000000000000000000110;
    n1464[914] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[913] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[912] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[911] = 42'b100000000000000000000010000000000000000000;
    n1464[910] = 42'b100000000000000000000010010000000000000000;
    n1464[909] = 42'b100000000000000000000010000010000000000000;
    n1464[908] = 42'b000000000000000000000000000000000000000000;
    n1464[907] = 42'b100100000000000000000000000000000000000110;
    n1464[906] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[905] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[904] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[903] = 42'b100000000000000000000010000000000000000000;
    n1464[902] = 42'b100000000000000000000010010000000000000000;
    n1464[901] = 42'b000000000000000000000000000000000000000000;
    n1464[900] = 42'b000000000000000000000000000000000000000000;
    n1464[899] = 42'b100000000000000000000000000000000000001100;
    n1464[898] = 42'b100000000000000000000010010000000000000010;
    n1464[897] = 42'b000000000000000000001000000000000000000000;
    n1464[896] = 42'b000000000000000000000000000000000000000010;
    n1464[895] = 42'b100000000000000000000010000000000000000000;
    n1464[894] = 42'b100000000000000000000010010000000000000010;
    n1464[893] = 42'b100000000000000000000000000000000000000000;
    n1464[892] = 42'b000000000000000000001000000000000000000010;
    n1464[891] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[890] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[889] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[888] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[887] = 42'b100000000000000000000010000000000000000000;
    n1464[886] = 42'b100000000000000000000010010000000000000000;
    n1464[885] = 42'b000000000000000000000000000000000000000000;
    n1464[884] = 42'b100000000000000000000000100000000000001100;
    n1464[883] = 42'b100000000000000000000001100010000000001100;
    n1464[882] = 42'b000000000000000000000000000110000000000000;
    n1464[881] = 42'b100010000000000000000000000000000000000110;
    n1464[880] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[879] = 42'b100000000000000000000010000000000000000000;
    n1464[878] = 42'b100000000000000000000010010000000000000000;
    n1464[877] = 42'b000000000000000000000000000000000000000000;
    n1464[876] = 42'b100000000000000000000000100000000000001100;
    n1464[875] = 42'b100000000000000000000001010010000000001100;
    n1464[874] = 42'b000000000000000000000000000000000000000000;
    n1464[873] = 42'b100010000000000000000000000000000000000110;
    n1464[872] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[871] = 42'b100000000000000000000010000000000000000000;
    n1464[870] = 42'b100000000000000000000010000000010000000000;
    n1464[869] = 42'b100000000000000000000010010000000000000000;
    n1464[868] = 42'b100000000000000000000010000010000000000000;
    n1464[867] = 42'b000000000000000000000000000000000000000000;
    n1464[866] = 42'b000000000000000000000000000000000000000000;
    n1464[865] = 42'b000000000000000000000000000000000000000000;
    n1464[864] = 42'b100000110001010000000000000000001010000110;
    n1464[863] = 42'b100000000000000000000010000000000000000000;
    n1464[862] = 42'b100000000000000000000010010000000000000000;
    n1464[861] = 42'b000000000000000000000000110000000000000000;
    n1464[860] = 42'b100110000000000000000000000000000000001110;
    n1464[859] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[858] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[857] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[856] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[855] = 42'b100000000000000000000010000000000000000000;
    n1464[854] = 42'b100000000000000000000010010000000000000000;
    n1464[853] = 42'b000000000000000000000000110000000000000000;
    n1464[852] = 42'b100010000000000000000000000000000000001110;
    n1464[851] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[850] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[849] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[848] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[847] = 42'b100000000000000000000010000000000000000000;
    n1464[846] = 42'b100000000000000000000010010000000000000000;
    n1464[845] = 42'b000000000000000000000001000000000000000000;
    n1464[844] = 42'b100100000000000000000000000000000000001110;
    n1464[843] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[842] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[841] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[840] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[839] = 42'b100000000000000000000010000000000000000000;
    n1464[838] = 42'b100000000000000000000010010000000000000000;
    n1464[837] = 42'b000000000000000000000000000000000000000000;
    n1464[836] = 42'b100000111011000000000000000000010000001100;
    n1464[835] = 42'b000000000000000000000000000000000000000000;
    n1464[834] = 42'b000000000000000000000000000000000000000000;
    n1464[833] = 42'b101000000000000000000000000000000000001110;
    n1464[832] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[831] = 42'b100000000000000000000010000000000000000000;
    n1464[830] = 42'b100000000000110010000000000000000010000010;
    n1464[829] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[828] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[827] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[826] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[825] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[824] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[823] = 42'b100000000000000000000010000000000000000000;
    n1464[822] = 42'b100000000000000000000010010000000000000000;
    n1464[821] = 42'b100000000000000000000011000010000000000000;
    n1464[820] = 42'b000000000000000000000000000110000000000000;
    n1464[819] = 42'b100010000000000000000000000000000000000110;
    n1464[818] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[817] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[816] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[815] = 42'b100000000000000000000010000000000000000000;
    n1464[814] = 42'b100000000000100000010000000000000000000010;
    n1464[813] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[812] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[811] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[810] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[809] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[808] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[807] = 42'b100000000000000000000010000000000000000000;
    n1464[806] = 42'b000000000000000000000000000000000000000010;
    n1464[805] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[804] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[803] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[802] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[801] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[800] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[799] = 42'b100000000000000000000010000000000000000000;
    n1464[798] = 42'b100000000000000000000010010000000000000000;
    n1464[797] = 42'b100000000000000000000010000010000000000000;
    n1464[796] = 42'b000000000000000000000000000000000000000000;
    n1464[795] = 42'b111110000000000000000000000000000000000110;
    n1464[794] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[793] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[792] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[791] = 42'b100000000000000000000010000000000000000000;
    n1464[790] = 42'b100000000000000000000010010000000000000000;
    n1464[789] = 42'b100000000000000000000010110010000000000000;
    n1464[788] = 42'b000000000000000000000000000110000000000000;
    n1464[787] = 42'b100010000000000000000000000000000000000110;
    n1464[786] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[785] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[784] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[783] = 42'b100000000000000000000010000000000000000000;
    n1464[782] = 42'b100000000000000000000010010000000000000000;
    n1464[781] = 42'b100000000000000000000010110010000000000000;
    n1464[780] = 42'b000000000000000000000000000110000000000000;
    n1464[779] = 42'b111110000000000000000000000000000000000110;
    n1464[778] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[777] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[776] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[775] = 42'b100000000000000000000010000000000000000000;
    n1464[774] = 42'b100000000000000000000010010000000000000000;
    n1464[773] = 42'b000000000000000000000000000000000000000000;
    n1464[772] = 42'b000000000000000000000000000000000000000000;
    n1464[771] = 42'b100000000000000000000000000000000000001100;
    n1464[770] = 42'b100000000000000000000010010000000000000010;
    n1464[769] = 42'b000000000000000000001000000000000000000000;
    n1464[768] = 42'b000000000000000000000000000000000000000010;
    n1464[767] = 42'b100000000000000000000010000000000000000000;
    n1464[766] = 42'b100000000000001000000010000000000010000010;
    n1464[765] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[764] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[763] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[762] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[761] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[760] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[759] = 42'b100000000000000000000010000000000000000000;
    n1464[758] = 42'b100000000000000000000010010000000000000000;
    n1464[757] = 42'b000000000000000000000000110000000000000000;
    n1464[756] = 42'b100000000000000000000000100000000000001100;
    n1464[755] = 42'b100000000000000000000001010010000000001100;
    n1464[754] = 42'b000000000000000000000000000000000000000000;
    n1464[753] = 42'b100000000000000010000000000000000010000110;
    n1464[752] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[751] = 42'b100000000000000000000010000000000000000000;
    n1464[750] = 42'b100000000000000100000010000000000010000010;
    n1464[749] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[748] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[747] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[746] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[745] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[744] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[743] = 42'b100000000000000000000010000000000000000000;
    n1464[742] = 42'b100000000000000000000010000000010000000000;
    n1464[741] = 42'b100000000000000000000010010000000000000000;
    n1464[740] = 42'b000000000000000000000000110000000000000000;
    n1464[739] = 42'b000000000000000000000000000000000000000000;
    n1464[738] = 42'b000000000000000000000000000000000000000000;
    n1464[737] = 42'b100000110001010000000000000000001010001110;
    n1464[736] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[735] = 42'b100000000000000000000010000000000000000000;
    n1464[734] = 42'b100000000000000000000010010000000000000000;
    n1464[733] = 42'b000000000000000000000000000000000000000000;
    n1464[732] = 42'b100000000000001000000000000000000010001110;
    n1464[731] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[730] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[729] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[728] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[727] = 42'b100000000000000000000010000000000000000000;
    n1464[726] = 42'b100000000000000000000010010000000000000000;
    n1464[725] = 42'b000000000000000000000000000000000000000000;
    n1464[724] = 42'b100000000000000010000000000000000010001110;
    n1464[723] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[722] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[721] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[720] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[719] = 42'b100000000000000000000010000000000000000000;
    n1464[718] = 42'b100000000000000000000010010000000000000000;
    n1464[717] = 42'b000000000000000000000000000000000000000000;
    n1464[716] = 42'b100000000000000100000000000000000010001110;
    n1464[715] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[714] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[713] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[712] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[711] = 42'b100000000000000000000010000000000000000000;
    n1464[710] = 42'b100000000000000000000010010000000000000000;
    n1464[709] = 42'b000000000000000000000000000000000000000000;
    n1464[708] = 42'b100000111011000000000000000000010000001100;
    n1464[707] = 42'b000000000000000000000000000000000000000000;
    n1464[706] = 42'b000000000000000000000000000000000000000000;
    n1464[705] = 42'b101000000000000000000000000000000000001110;
    n1464[704] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[703] = 42'b100000000000000000000010000000000000000000;
    n1464[702] = 42'b100000000000011000000000000000000010000010;
    n1464[701] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[700] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[699] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[698] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[697] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[696] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[695] = 42'b100000000000000000000010000000000000000000;
    n1464[694] = 42'b100000000000000010000010000000000010000010;
    n1464[693] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[692] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[691] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[690] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[689] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[688] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[687] = 42'b100000000000000000000010000000000000000000;
    n1464[686] = 42'b100000000000010100000000000000000010000010;
    n1464[685] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[684] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[683] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[682] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[681] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[680] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[679] = 42'b100000000000000000000010000000000000000000;
    n1464[678] = 42'b000000000000000000000000000000000000000010;
    n1464[677] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[676] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[675] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[674] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[673] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[672] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[671] = 42'b100000000000000000000010000000000000000000;
    n1464[670] = 42'b100000000000000000000010010000000000000000;
    n1464[669] = 42'b100000000000000000000010000010000000000000;
    n1464[668] = 42'b000000000000000000000000000000000000000000;
    n1464[667] = 42'b100000000000001000000000000000000010000110;
    n1464[666] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[665] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[664] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[663] = 42'b100000000000000000000010000000000000000000;
    n1464[662] = 42'b100000000000000000000010010000000000000000;
    n1464[661] = 42'b100000000000000000000010000010000000000000;
    n1464[660] = 42'b000000000000000000000000000000000000000000;
    n1464[659] = 42'b100000000000000010000000000000000010000110;
    n1464[658] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[657] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[656] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[655] = 42'b100000000000000000000010000000000000000000;
    n1464[654] = 42'b100000000000000000000010010000000000000000;
    n1464[653] = 42'b100000000000000000000010000010000000000000;
    n1464[652] = 42'b000000000000000000000000000000000000000000;
    n1464[651] = 42'b100000000000000100000000000000000010000110;
    n1464[650] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[649] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[648] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[647] = 42'b100000000000000000000010000000000000000000;
    n1464[646] = 42'b100000000000000000000010010000000000000000;
    n1464[645] = 42'b000000000000000000000000000000000000000000;
    n1464[644] = 42'b000000000000000000000000000000000000000000;
    n1464[643] = 42'b100000000000000000000000000000000000001100;
    n1464[642] = 42'b100000000000000000000010010000000000000010;
    n1464[641] = 42'b000000000000000000001000000000000000000000;
    n1464[640] = 42'b000000000000000000000000000000000000000010;
    n1464[639] = 42'b100000000000000000000010000000000000000000;
    n1464[638] = 42'b100000000000000000000010010000000000000010;
    n1464[637] = 42'b100000000000000000000000000000000000000000;
    n1464[636] = 42'b000000000000000000001000000000000000000010;
    n1464[635] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[634] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[633] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[632] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[631] = 42'b100000000000000000000010000000000000000000;
    n1464[630] = 42'b100000000000000000000010010000000000000000;
    n1464[629] = 42'b000000000000000000000000000000000000000000;
    n1464[628] = 42'b100000000000000000000000100000000000001100;
    n1464[627] = 42'b100000000000000000000001100010000000001100;
    n1464[626] = 42'b000000000000000000000000000110000000000000;
    n1464[625] = 42'b100000000000000010000000000000000010000110;
    n1464[624] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[623] = 42'b100000000000000000000010000000000000000000;
    n1464[622] = 42'b100000000000000000000010010000000000000000;
    n1464[621] = 42'b000000000000000000000000000000000000000000;
    n1464[620] = 42'b100000000000000000000000100000000000001100;
    n1464[619] = 42'b100000000000000000000001010010000000001100;
    n1464[618] = 42'b000000000000000000000000000000000000000000;
    n1464[617] = 42'b100000000000000010000000000000000010000110;
    n1464[616] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[615] = 42'b100000000000000000000010000000000000000000;
    n1464[614] = 42'b100000000000000000000010000000010000000000;
    n1464[613] = 42'b100000000000000000000010010000000000000000;
    n1464[612] = 42'b100000000000000000000010110010000000000000;
    n1464[611] = 42'b000000000000000000000000000110000000000000;
    n1464[610] = 42'b000000000000000000000000000000000000000000;
    n1464[609] = 42'b000000000000000000000000000000000000000000;
    n1464[608] = 42'b100000110001010000000000000000001010000110;
    n1464[607] = 42'b100000000000000000000010000000000000000000;
    n1464[606] = 42'b100000000000000000000010010000000000000000;
    n1464[605] = 42'b000000000000000000000000110000000000000000;
    n1464[604] = 42'b100000000000001000000000000000000010001110;
    n1464[603] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[602] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[601] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[600] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[599] = 42'b100000000000000000000010000000000000000000;
    n1464[598] = 42'b100000000000000000000010010000000000000000;
    n1464[597] = 42'b000000000000000000000000110000000000000000;
    n1464[596] = 42'b100000000000000010000000000000000010001110;
    n1464[595] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[594] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[593] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[592] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[591] = 42'b100000000000000000000010000000000000000000;
    n1464[590] = 42'b100000000000000000000010010000000000000000;
    n1464[589] = 42'b000000000000000000000001000000000000000000;
    n1464[588] = 42'b100000000000000100000000000000000010001110;
    n1464[587] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[586] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[585] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[584] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[583] = 42'b100000000000000000000010000000000000000000;
    n1464[582] = 42'b100000000000000000000010010000000000000000;
    n1464[581] = 42'b000000000000000000000000000000000000000000;
    n1464[580] = 42'b100000111011000000000000000000010000001100;
    n1464[579] = 42'b000000000000000000000000000000000000000000;
    n1464[578] = 42'b000000000000000000000000000000000000000000;
    n1464[577] = 42'b101000000000000000000000000000000000001110;
    n1464[576] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[575] = 42'b100000000000000000000010000000000000000000;
    n1464[574] = 42'b100000000000000000000000000000001000000010;
    n1464[573] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[572] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[571] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[570] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[569] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[568] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[567] = 42'b100000000000000000000010000000000000000000;
    n1464[566] = 42'b100000000000000000000010010000000000000000;
    n1464[565] = 42'b100000000000000000000011000010000000000000;
    n1464[564] = 42'b000000000000000000000000000110000000000000;
    n1464[563] = 42'b100000000000000010000000000000000010000110;
    n1464[562] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[561] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[560] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[559] = 42'b100000000000000000000010000000000000000000;
    n1464[558] = 42'b100000000001000100000000000000000010000010;
    n1464[557] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[556] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[555] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[554] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[553] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[552] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[551] = 42'b100000000000000000000010000000000000000000;
    n1464[550] = 42'b000000000000000000000000000000000000000010;
    n1464[549] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[548] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[547] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[546] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[545] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[544] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[543] = 42'b100000000000000000000010000000000000000000;
    n1464[542] = 42'b100000000000000000000010010000000000000000;
    n1464[541] = 42'b100000000000000000000010110010000000000000;
    n1464[540] = 42'b000000000000000000000000000110000000000000;
    n1464[539] = 42'b100000000000001000000000000000000010000110;
    n1464[538] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[537] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[536] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[535] = 42'b100000000000000000000010000000000000000000;
    n1464[534] = 42'b100000000000000000000010010000000000000000;
    n1464[533] = 42'b100000000000000000000010110010000000000000;
    n1464[532] = 42'b000000000000000000000000000110000000000000;
    n1464[531] = 42'b100000000000000010000000000000000010000110;
    n1464[530] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[529] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[528] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[527] = 42'b100000000000000000000010000000000000000000;
    n1464[526] = 42'b100000000000000000000010010000000000000000;
    n1464[525] = 42'b100000000000000000000011000010000000000000;
    n1464[524] = 42'b000000000000000000000000000110000000000000;
    n1464[523] = 42'b100000000000000100000000000000000010000110;
    n1464[522] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[521] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[520] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[519] = 42'b100000000000000000000010000000000000000000;
    n1464[518] = 42'b100000000000000000000010010000000000000000;
    n1464[517] = 42'b000000000000000000000000000000000000000000;
    n1464[516] = 42'b000000000000000000000000000000000000000000;
    n1464[515] = 42'b100000000000000000000000000000000000001100;
    n1464[514] = 42'b100000000000000000000010010000000000000010;
    n1464[513] = 42'b000000000000000000001000000000000000000000;
    n1464[512] = 42'b000000000000000000000000000000000000000010;
    n1464[511] = 42'b100000000000000000000010000000000000000000;
    n1464[510] = 42'b100000111100110000000010000000001010000010;
    n1464[509] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[508] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[507] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[506] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[505] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[504] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[503] = 42'b100000000000000000000010000000000000000000;
    n1464[502] = 42'b100000000000000000000010010000000000000000;
    n1464[501] = 42'b000000000000000000000000110000000000000000;
    n1464[500] = 42'b100000000000000000000000100000000000001100;
    n1464[499] = 42'b100000000000000000000001010010000000001100;
    n1464[498] = 42'b000000000000000000000000000000000000000000;
    n1464[497] = 42'b100000111100010000000000000000001010000110;
    n1464[496] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[495] = 42'b100000000000000000000010000000000000000000;
    n1464[494] = 42'b100000000011111000000000000000000000000010;
    n1464[493] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[492] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[491] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[490] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[489] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[488] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[487] = 42'b100000000000000000000010000000000000000000;
    n1464[486] = 42'b100110000000000000110000000000000000001000;
    n1464[485] = 42'b100010000000000000110000000000000000001000;
    n1464[484] = 42'b100100000000000000000000000000000000001000;
    n1464[483] = 42'b100000000000000100000010000000000000000000;
    n1464[482] = 42'b100000000000000000000010000000000000100000;
    n1464[481] = 42'b100000000000001000000010000000000000000000;
    n1464[480] = 42'b100000000000000000000010000000000001000000;
    n1464[479] = 42'b100000000000000000000010000000000000000000;
    n1464[478] = 42'b100000000000000000000010010000000000000000;
    n1464[477] = 42'b000000000000000000000000000000000000000000;
    n1464[476] = 42'b100000111100110000000000000000001010001110;
    n1464[475] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[474] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[473] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[472] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[471] = 42'b100000000000000000000010000000000000000000;
    n1464[470] = 42'b100000000000000000000010010000000000000000;
    n1464[469] = 42'b000000000000000000000000000000000000000000;
    n1464[468] = 42'b100000111100010000000000000000001010001110;
    n1464[467] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[466] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[465] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[464] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[463] = 42'b100000000000000000000010000000000000000000;
    n1464[462] = 42'b100000000000000000000010010000000000000000;
    n1464[461] = 42'b000000000000000000000000000000000000000000;
    n1464[460] = 42'b100000011000000000000000000000010010001100;
    n1464[459] = 42'b000000000000000000000000000000000000000000;
    n1464[458] = 42'b101000000000000000000000000000000000001110;
    n1464[457] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[456] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[455] = 42'b100000000000000000000010000000000000000000;
    n1464[454] = 42'b100000000000000000000010010000000000000000;
    n1464[453] = 42'b000000000000000000000000000000000000000000;
    n1464[452] = 42'b100000111011000000000000000000010000001100;
    n1464[451] = 42'b000000000000000000000000000000000000000000;
    n1464[450] = 42'b000000000000000000000000000000000000000000;
    n1464[449] = 42'b101000000000000000000000000000000000001110;
    n1464[448] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[447] = 42'b100000000000000000000010000000000000000000;
    n1464[446] = 42'b100000011100111000000000000000000010000010;
    n1464[445] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[444] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[443] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[442] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[441] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[440] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[439] = 42'b100000000000000000000010000000000000000000;
    n1464[438] = 42'b100000111100010000000010000000001010000010;
    n1464[437] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[436] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[435] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[434] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[433] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[432] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[431] = 42'b100000000000000000000010000000000000000000;
    n1464[430] = 42'b100000011000100100000000000000000010000010;
    n1464[429] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[428] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[427] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[426] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[425] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[424] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[423] = 42'b100000000000000000000010000000000000000000;
    n1464[422] = 42'b000000000000000000000000000000000000000010;
    n1464[421] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[420] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[419] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[418] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[417] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[416] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[415] = 42'b100000000000000000000010000000000000000000;
    n1464[414] = 42'b100000000000000000000010010000000000000000;
    n1464[413] = 42'b100000000000000000000010000010000000000000;
    n1464[412] = 42'b000000000000000000000000000000000000000000;
    n1464[411] = 42'b100000111100110000000000000000001010000110;
    n1464[410] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[409] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[408] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[407] = 42'b100000000000000000000010000000000000000000;
    n1464[406] = 42'b100000000000000000000010010000000000000000;
    n1464[405] = 42'b100000000000000000000010000010000000000000;
    n1464[404] = 42'b000000000000000000000000000000000000000000;
    n1464[403] = 42'b100000111100010000000000000000001010000110;
    n1464[402] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[401] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[400] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[399] = 42'b100000000000000000000010000000000000000000;
    n1464[398] = 42'b100000000000000000000010010000000000000000;
    n1464[397] = 42'b100000000000000000000010000010000000000000;
    n1464[396] = 42'b000000000000000000000000000000000000000000;
    n1464[395] = 42'b100000011000000000000000000000010010000100;
    n1464[394] = 42'b000000000000000000000000000000000000000000;
    n1464[393] = 42'b101000000000000000000000000000000000000110;
    n1464[392] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[391] = 42'b100000000000000000000010000000000000000000;
    n1464[390] = 42'b100000000000000000000010010000000000000000;
    n1464[389] = 42'b000000000000000000000000000000000000000000;
    n1464[388] = 42'b000000000000000000000000000000000000000000;
    n1464[387] = 42'b100000000000000000000000000000000000001100;
    n1464[386] = 42'b100000000000000000000010010000000000000010;
    n1464[385] = 42'b000000000000000000001000000000000000000000;
    n1464[384] = 42'b000000000000000000000000000000000000000010;
    n1464[383] = 42'b100000000000000000000010000000000000000000;
    n1464[382] = 42'b100000000000000000000010010000000000000010;
    n1464[381] = 42'b000000000000000000000000000000000000000000;
    n1464[380] = 42'b000000000000000000001000000000000000000010;
    n1464[379] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[378] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[377] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[376] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[375] = 42'b100000000000000000000010000000000000000000;
    n1464[374] = 42'b100000000000000000000010010000000000000000;
    n1464[373] = 42'b000000000000000000000000000000000000000000;
    n1464[372] = 42'b100000000000000000000000100000000000001100;
    n1464[371] = 42'b100000000000000000000001100010000000001100;
    n1464[370] = 42'b000000000000000000000000000110000000000000;
    n1464[369] = 42'b100000111100010000000000000000001010000110;
    n1464[368] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[367] = 42'b100000000000000000000010000000000000000000;
    n1464[366] = 42'b100000000000000000000010010000000000000000;
    n1464[365] = 42'b000000000000000000000000000000000000000000;
    n1464[364] = 42'b100000000000000000000000100000000000001100;
    n1464[363] = 42'b100000000000000000000001010010000000001100;
    n1464[362] = 42'b000000000000000000000000000000000000000000;
    n1464[361] = 42'b100000111100010000000000000000001010000110;
    n1464[360] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[359] = 42'b100000000000000000000010000000000000000000;
    n1464[358] = 42'b100110000000000000110000000000000000001000;
    n1464[357] = 42'b100010000000000000110000000000000000001000;
    n1464[356] = 42'b100100000000000000000000000000000000001000;
    n1464[355] = 42'b100000000000000100000010000000000000000000;
    n1464[354] = 42'b100000000000000000000010000000000000100000;
    n1464[353] = 42'b100000000000001000000010000000000000000000;
    n1464[352] = 42'b100000000000000000000010000000000001000000;
    n1464[351] = 42'b100000000000000000000010000000000000000000;
    n1464[350] = 42'b100000000000000000000000000000000000000000;
    n1464[349] = 42'b000000000000000000000000000000000000000010;
    n1464[348] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[347] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[346] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[345] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[344] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[343] = 42'b100000000000000000000010000000000000000000;
    n1464[342] = 42'b100000000000000000000010010000000000000000;
    n1464[341] = 42'b000000000000000000000000110000000000000000;
    n1464[340] = 42'b100000111100010000000000000000001010001110;
    n1464[339] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[338] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[337] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[336] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[335] = 42'b100000000000000000000010000000000000000000;
    n1464[334] = 42'b100000000000000000000010010000000000000000;
    n1464[333] = 42'b000000000000000000000000110000000000000000;
    n1464[332] = 42'b100000011000000000000000000000010010001100;
    n1464[331] = 42'b000000000000000000000000000000000000000000;
    n1464[330] = 42'b101000000000000000000000000000000000001110;
    n1464[329] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[328] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[327] = 42'b100000000000000000000010000000000000000000;
    n1464[326] = 42'b100000000000000000000010010000000000000000;
    n1464[325] = 42'b000000000000000000000000000000000000000000;
    n1464[324] = 42'b100000111011000000000000000000010000001100;
    n1464[323] = 42'b000000000000000000000000000000000000000000;
    n1464[322] = 42'b000000000000000000000000000000000000000000;
    n1464[321] = 42'b101000000000000000000000000000000000001110;
    n1464[320] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[319] = 42'b100000000000000000000010000000000000000000;
    n1464[318] = 42'b100000000000000000000000000000001000000010;
    n1464[317] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[316] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[315] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[314] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[313] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[312] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[311] = 42'b100000000000000000000010000000000000000000;
    n1464[310] = 42'b100000000000000000000010010000000000000000;
    n1464[309] = 42'b100000000000000000000011000010000000000000;
    n1464[308] = 42'b000000000000000000000000000110000000000000;
    n1464[307] = 42'b100000111100010000000000000000001010000110;
    n1464[306] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[305] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[304] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[303] = 42'b100000000000000000000010000000000000000000;
    n1464[302] = 42'b100000000000000000000000000000000000000000;
    n1464[301] = 42'b100100000000000000110000000000000000001010;
    n1464[300] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[299] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[298] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[297] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[296] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[295] = 42'b100000000000000000000010000000000000000000;
    n1464[294] = 42'b000000000000000000000000000000000000000010;
    n1464[293] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[292] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[291] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[290] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[289] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[288] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[287] = 42'b100000000000000000000010000000000000000000;
    n1464[286] = 42'b000000000000000000000000000000000000000010;
    n1464[285] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[284] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[283] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[282] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[281] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[280] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[279] = 42'b100000000000000000000010000000000000000000;
    n1464[278] = 42'b100000000000000000000010010000000000000000;
    n1464[277] = 42'b100000000000000000000010110010000000000000;
    n1464[276] = 42'b000000000000000000000000000110000000000000;
    n1464[275] = 42'b100000111100010000000000000000001010000110;
    n1464[274] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[273] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[272] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[271] = 42'b100000000000000000000010000000000000000000;
    n1464[270] = 42'b100000000000000000000010010000000000000000;
    n1464[269] = 42'b100000000000000000000010110010000000000000;
    n1464[268] = 42'b000000000000000000000000000110000000000000;
    n1464[267] = 42'b100000011000000000000000000000010010000100;
    n1464[266] = 42'b000000000000000000000000000000000000000000;
    n1464[265] = 42'b101000000000000000000000000000000000000110;
    n1464[264] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[263] = 42'b100000000000000000000010000000000000000000;
    n1464[262] = 42'b100000000000000000000010010000000000000000;
    n1464[261] = 42'b000000000000000000000000000000000000000000;
    n1464[260] = 42'b000000000000000000000000000000000000000000;
    n1464[259] = 42'b100000000000000000000000000000000000001100;
    n1464[258] = 42'b100000000000000000000010010000000000000010;
    n1464[257] = 42'b000000000000000000001000000000000000000000;
    n1464[256] = 42'b000000000000000000000000000000000000000010;
    n1464[255] = 42'b100000000000000000000010000000000000000000;
    n1464[254] = 42'b100000111100100000000010000000001010000010;
    n1464[253] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[252] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[251] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[250] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[249] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[248] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[247] = 42'b100000000000000000000010000000000000000000;
    n1464[246] = 42'b100000000000000000000010010000000000000000;
    n1464[245] = 42'b000000000000000000000000110000000000000000;
    n1464[244] = 42'b100000000000000000000000100000000000001100;
    n1464[243] = 42'b100000000000000000000001010010000000001100;
    n1464[242] = 42'b000000000000000000000000000000000000000000;
    n1464[241] = 42'b100000010100010010000000000000001010000101;
    n1464[240] = 42'b000000000000000000000000000000000000000010;
    n1464[239] = 42'b100000000000000000000010000000000000000000;
    n1464[238] = 42'b000000000000000000000000000000000000000010;
    n1464[237] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[236] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[235] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[234] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[233] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[232] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[231] = 42'b100000000000000000000010000000000000000000;
    n1464[230] = 42'b100110000000000000110000000000000000001000;
    n1464[229] = 42'b100010000000000000110000000000000000001000;
    n1464[228] = 42'b100100000000000000000000000000000000001000;
    n1464[227] = 42'b100000000000000100000010000000000000000000;
    n1464[226] = 42'b100000000000000000000010000000000000100000;
    n1464[225] = 42'b100000000000001000000010000000000000000000;
    n1464[224] = 42'b100000000000000000000010000000000001000000;
    n1464[223] = 42'b100000000000000000000010000000000000000000;
    n1464[222] = 42'b100000000000000000000010010000000000000000;
    n1464[221] = 42'b000000000000000000000000000000000000000000;
    n1464[220] = 42'b100000111100100000000000000000001010001110;
    n1464[219] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[218] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[217] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[216] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[215] = 42'b100000000000000000000010000000000000000000;
    n1464[214] = 42'b100000000000000000000010010000000000000000;
    n1464[213] = 42'b000000000000000000000000000000000000000000;
    n1464[212] = 42'b100000010100010010000000000000001010001101;
    n1464[211] = 42'b000000000000000000000000000000000000000010;
    n1464[210] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[209] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[208] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[207] = 42'b100000000000000000000010000000000000000000;
    n1464[206] = 42'b100000000000000000000010010000000000000000;
    n1464[205] = 42'b000000000000000000000000000000000000000000;
    n1464[204] = 42'b100000011100000000000000000000010010001100;
    n1464[203] = 42'b000000000000000000000000000000000000000000;
    n1464[202] = 42'b101000000000000000000000000000000000001110;
    n1464[201] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[200] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[199] = 42'b100000000000000000000010000000000000000000;
    n1464[198] = 42'b100000000000000000000010010000000000000000;
    n1464[197] = 42'b000000000000000000000000000000000000000000;
    n1464[196] = 42'b100000111011000000000000000000010000001100;
    n1464[195] = 42'b000000000000000000000000000000000000000000;
    n1464[194] = 42'b000000000000000000000000000000000000000000;
    n1464[193] = 42'b101000000000000000000000000000000000001110;
    n1464[192] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[191] = 42'b100000000000000000000010000000000000000000;
    n1464[190] = 42'b100000011100100100000000000000000010000010;
    n1464[189] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[188] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[187] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[186] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[185] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[184] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[183] = 42'b100000000000000000000010000000000000000000;
    n1464[182] = 42'b100000010100010010000010000000001010000001;
    n1464[181] = 42'b000000000000000000000000000000000000000010;
    n1464[180] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[179] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[178] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[177] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[176] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[175] = 42'b100000000000000000000010000000000000000000;
    n1464[174] = 42'b100000000000000000000000000000000000000010;
    n1464[173] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[172] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[171] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[170] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[169] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[168] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[167] = 42'b100000000000000000000010000000000000000000;
    n1464[166] = 42'b000000000000000000000000000000000000000010;
    n1464[165] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[164] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[163] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[162] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[161] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[160] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[159] = 42'b100000000000000000000010000000000000000000;
    n1464[158] = 42'b100000000000000000000010010000000000000000;
    n1464[157] = 42'b100000000000000000000010000010000000000000;
    n1464[156] = 42'b000000000000000000000000000000000000000000;
    n1464[155] = 42'b100000111100100000000000000000001010000110;
    n1464[154] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[153] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[152] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[151] = 42'b100000000000000000000010000000000000000000;
    n1464[150] = 42'b100000000000000000000010010000000000000000;
    n1464[149] = 42'b100000000000000000000010000010000000000000;
    n1464[148] = 42'b000000000000000000000000000000000000000000;
    n1464[147] = 42'b100000010100010010000000000000001010000110;
    n1464[146] = 42'b000000000000000000000000000000000000000010;
    n1464[145] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[144] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[143] = 42'b100000000000000000000010000000000000000000;
    n1464[142] = 42'b100000000000000000000010010000000000000000;
    n1464[141] = 42'b100000000000000000000010000010000000000000;
    n1464[140] = 42'b000000000000000000000000000000000000000000;
    n1464[139] = 42'b100000011100000000000000000000010010000100;
    n1464[138] = 42'b000000000000000000000000000000000000000000;
    n1464[137] = 42'b101000000000000000000000000000000000000110;
    n1464[136] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[135] = 42'b100000000000000000000010000000000000000000;
    n1464[134] = 42'b100000000000000000000010010000000000000000;
    n1464[133] = 42'b000000000000000000000000000000000000000000;
    n1464[132] = 42'b000000000000000000000000000000000000000000;
    n1464[131] = 42'b100000000000000000000000000000000000001100;
    n1464[130] = 42'b100000000000000000000010010000000000000010;
    n1464[129] = 42'b000000000000000000001000000000000000000000;
    n1464[128] = 42'b000000000000000000000000000000000000000010;
    n1464[127] = 42'b100000000000000000000010000000000000000000;
    n1464[126] = 42'b100000000000000000000010010000000000000010;
    n1464[125] = 42'b100000000000000000000000000000000000000000;
    n1464[124] = 42'b000000000000000000001000000000000000000010;
    n1464[123] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[122] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[121] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[120] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[119] = 42'b100000000000000000000010000000000000000000;
    n1464[118] = 42'b100000000000000000000010010000000000000000;
    n1464[117] = 42'b000000000000000000000000000000000000000000;
    n1464[116] = 42'b100000000000000000000000100000000000001100;
    n1464[115] = 42'b100000000000000000000001100010000000001100;
    n1464[114] = 42'b000000000000000000000000000110000000000000;
    n1464[113] = 42'b100000010100010010000000000000001010000101;
    n1464[112] = 42'b000000000000000000000000000000000000000010;
    n1464[111] = 42'b100000000000000000000010000000000000000000;
    n1464[110] = 42'b100000000000000000000010010000000000000000;
    n1464[109] = 42'b000000000000000000000000000000000000000000;
    n1464[108] = 42'b100000000000000000000000100000000000001100;
    n1464[107] = 42'b100000000000000000000001010010000000001100;
    n1464[106] = 42'b000000000000000000000000000000000000000000;
    n1464[105] = 42'b100000010100010010000000000000001010000101;
    n1464[104] = 42'b000000000000000000000000000000000000000010;
    n1464[103] = 42'b100000000000000000000010000000000000000000;
    n1464[102] = 42'b100110000000000000110000000000000000001000;
    n1464[101] = 42'b100010000000000000110000000000000000001000;
    n1464[100] = 42'b100100000000000000000000000000000000001000;
    n1464[99] = 42'b100000000000000100000010000000000000000000;
    n1464[98] = 42'b100000000000000000000010000000000000100000;
    n1464[97] = 42'b100000000000001000000010000000000000000000;
    n1464[96] = 42'b100000000000000000000010000000000001000000;
    n1464[95] = 42'b100000000000000000000010000000000000000000;
    n1464[94] = 42'b100000000000000000000000000000001100000010;
    n1464[93] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[92] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[91] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[90] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[89] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[88] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[87] = 42'b100000000000000000000010000000000000000000;
    n1464[86] = 42'b100000000000000000000010010000000000000000;
    n1464[85] = 42'b000000000000000000000000110000000000000000;
    n1464[84] = 42'b100000010100010010000000000000001010001101;
    n1464[83] = 42'b000000000000000000000000000000000000000010;
    n1464[82] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[81] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[80] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[79] = 42'b100000000000000000000010000000000000000000;
    n1464[78] = 42'b100000000000000000000010010000000000000000;
    n1464[77] = 42'b000000000000000000000000110000000000000000;
    n1464[76] = 42'b100000011100000000000000000000010010001100;
    n1464[75] = 42'b000000000000000000000000000000000000000000;
    n1464[74] = 42'b101000000000000000000000000000000000001110;
    n1464[73] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[72] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[71] = 42'b100000000000000000000010000000000000000000;
    n1464[70] = 42'b100000000000000000000010010000000000000000;
    n1464[69] = 42'b000000000000000000000000000000000000000000;
    n1464[68] = 42'b100000111011000000000000000000010000001100;
    n1464[67] = 42'b000000000000000000000000000000000000000000;
    n1464[66] = 42'b000000000000000000000000000000000000000000;
    n1464[65] = 42'b101000000000000000000000000000000000001110;
    n1464[64] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[63] = 42'b100000000000000000000010000000000000000000;
    n1464[62] = 42'b100000000000000000000000000000001000000010;
    n1464[61] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[60] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[59] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[58] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[57] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[56] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[55] = 42'b100000000000000000000010000000000000000000;
    n1464[54] = 42'b100000000000000000000010010000000000000000;
    n1464[53] = 42'b100000000000000000000011000010000000000000;
    n1464[52] = 42'b000000000000000000000000000110000000000000;
    n1464[51] = 42'b100000010100010010000000000000001010000101;
    n1464[50] = 42'b000000000000000000000000000000000000000010;
    n1464[49] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[48] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[47] = 42'b100000000000000000000010000000000000000000;
    n1464[46] = 42'b000000000000000000000000000000000000000000;
    n1464[45] = 42'b000000000000000000100000000000000000000000;
    n1464[44] = 42'b100000000000000100000000000000000010001010;
    n1464[43] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[42] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[41] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[40] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[39] = 42'b100000000000000000000010000000000000000000;
    n1464[38] = 42'b000000000000000000000000000000000000000010;
    n1464[37] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[36] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[35] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[34] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[33] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[32] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[31] = 42'b100000000000000000000010000000000000000000;
    n1464[30] = 42'b000000000000000000000000000000000000000010;
    n1464[29] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[28] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[27] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[26] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[25] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[24] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[23] = 42'b100000000000000000000010000000000000000000;
    n1464[22] = 42'b100000000000000000000010010000000000000000;
    n1464[21] = 42'b100000000000000000000010110010000000000000;
    n1464[20] = 42'b000000000000000000000000000110000000000000;
    n1464[19] = 42'b100000010100010010000000000000001010000101;
    n1464[18] = 42'b000000000000000000000000000000000000000010;
    n1464[17] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[16] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[15] = 42'b100000000000000000000010000000000000000000;
    n1464[14] = 42'b100000000000000000000010010000000000000000;
    n1464[13] = 42'b100000000000000000000010110010000000000000;
    n1464[12] = 42'b000000000000000000000000000110000000000000;
    n1464[11] = 42'b100000011100000000000000000000010010000100;
    n1464[10] = 42'b000000000000000000000000000000000000000000;
    n1464[9] = 42'b101000000000000000000000000000000000000110;
    n1464[8] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1464[7] = 42'b100000000000000000000010000000000000000000;
    n1464[6] = 42'b100000000000000000000010010000000000000000;
    n1464[5] = 42'b000000000000000000000000000000000000000000;
    n1464[4] = 42'b000000000000000000000000000000000000000000;
    n1464[3] = 42'b100000000000000000000000000000000000001100;
    n1464[2] = 42'b100000000000000000000010010000000000000010;
    n1464[1] = 42'b000000000000000000001000000000000000000000;
    n1464[0] = 42'b000000000000000000000000000000000000000010;
    end
  assign n1465_data = n1464[n1405_o];
  /* HUC6280_MC.vhd:6984:54  */
  /* HUC6280_MC.vhd:6984:53  */
  reg [41:0] n1466[2047:0] ; // memory
  initial begin
    n1466[2047] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2046] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2045] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2044] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2043] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2042] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2041] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2040] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2039] = 42'b100000000000000000000010010000000000000000;
    n1466[2038] = 42'b000000000000000000000000110000000000000000;
    n1466[2037] = 42'b100000000000000000000000100000000000001100;
    n1466[2036] = 42'b100000000000000000000001010010000000001100;
    n1466[2035] = 42'b000000000000000000000000000000000000000000;
    n1466[2034] = 42'b100000000000000000000000000000010000000100;
    n1466[2033] = 42'b000000000000000000000001110000000000000000;
    n1466[2032] = 42'b100000001001010000000000000000010010001100;
    n1466[2031] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2030] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2029] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2028] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2027] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2026] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2025] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2024] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2023] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2022] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2021] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2020] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2019] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2018] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2017] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2016] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2015] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2014] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2013] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2012] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2011] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2010] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2009] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2008] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2007] = 42'b100000000000000000000010010000000000000000;
    n1466[2006] = 42'b000000000000000000000000000000000000000000;
    n1466[2005] = 42'b100000000000000000000000000000010000001100;
    n1466[2004] = 42'b000000000000000000000001110000000000000000;
    n1466[2003] = 42'b100000001001010000000000000000010010001100;
    n1466[2002] = 42'b101000000000000000000000000000000000001110;
    n1466[2001] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2000] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1999] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1998] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1997] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1996] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1995] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1994] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1993] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1992] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1991] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1990] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1989] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1988] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1987] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1986] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1985] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1984] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1983] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1982] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1981] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1980] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1979] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1978] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1977] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1976] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1975] = 42'b100000000000000000000010000000010000000000;
    n1466[1974] = 42'b000000000000000000000001110000000000000000;
    n1466[1973] = 42'b100000001001010000000000000000010010001100;
    n1466[1972] = 42'b101000000000000000000000000000000000001110;
    n1466[1971] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1970] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1969] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1968] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1967] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1966] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1965] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1964] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1963] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1962] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1961] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1960] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1959] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1958] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1957] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1956] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1955] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1954] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1953] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1952] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1951] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1950] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1949] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1948] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1947] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1946] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1945] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1944] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1943] = 42'b100000000000000000000010010000000000000000;
    n1466[1942] = 42'b100000000000000000000010000010000000000000;
    n1466[1941] = 42'b000000000000000000000000000000000000000000;
    n1466[1940] = 42'b100000000000000000000000000000010000000100;
    n1466[1939] = 42'b000000000000000000000001110000000000000000;
    n1466[1938] = 42'b100000001001010000000000000000010010001100;
    n1466[1937] = 42'b101000000000000000000000000000000000001110;
    n1466[1936] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1935] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1934] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1933] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1932] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1931] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1930] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1929] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1928] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1927] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1926] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1925] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1924] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1923] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1922] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1921] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1920] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1919] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1918] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1917] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1916] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1915] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1914] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1913] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1912] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1911] = 42'b100000000000000000000010010000000000000000;
    n1466[1910] = 42'b000000000000000000000000000000000000000000;
    n1466[1909] = 42'b100000000000000000000000100000000000001100;
    n1466[1908] = 42'b100000000000000000000001100010000000001100;
    n1466[1907] = 42'b000000000000000000000000000110000000000000;
    n1466[1906] = 42'b100000000000000000000000000000010000000100;
    n1466[1905] = 42'b000000000000000000000001110000000000000000;
    n1466[1904] = 42'b100000001001010000000000000000010010001100;
    n1466[1903] = 42'b100000000000000000000010010000000000000000;
    n1466[1902] = 42'b000000000000000000000000000000000000000000;
    n1466[1901] = 42'b100000000000000000000000100000000000001100;
    n1466[1900] = 42'b100000000000000000000001010010000000001100;
    n1466[1899] = 42'b000000000000000000000000000000000000000000;
    n1466[1898] = 42'b100000000000000000000000000000010000000100;
    n1466[1897] = 42'b000000000000000000000001110000000000000000;
    n1466[1896] = 42'b100000001001010000000000000000010010001100;
    n1466[1895] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1894] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1893] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1892] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1891] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1890] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1889] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1888] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1887] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1886] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1885] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1884] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1883] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1882] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1881] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1880] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1879] = 42'b100000000000000000000010010000000000000000;
    n1466[1878] = 42'b000000000000000000000000110000000000000000;
    n1466[1877] = 42'b100000000000000000000000000000010000001100;
    n1466[1876] = 42'b000000000000000000000001110000000000000000;
    n1466[1875] = 42'b100000001001010000000000000000010010001100;
    n1466[1874] = 42'b101000000000000000000000000000000000001110;
    n1466[1873] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1872] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1871] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1870] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1869] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1868] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1867] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1866] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1865] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1864] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1863] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1862] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1861] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1860] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1859] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1858] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1857] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1856] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1855] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1854] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1853] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1852] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1851] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1850] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1849] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1848] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1847] = 42'b100000000000000000000010010000000000000000;
    n1466[1846] = 42'b100000000000000000000011000010000000000000;
    n1466[1845] = 42'b000000000000000000000000000110000000000000;
    n1466[1844] = 42'b100000000000000000000000000000010000000100;
    n1466[1843] = 42'b000000000000000000000001110000000000000000;
    n1466[1842] = 42'b100000001001010000000000000000010010001100;
    n1466[1841] = 42'b101000000000000000000000000000000000001110;
    n1466[1840] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1839] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1838] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1837] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1836] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1835] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1834] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1833] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1832] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1831] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1830] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1829] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1828] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1827] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1826] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1825] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1824] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1823] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1822] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1821] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1820] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1819] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1818] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1817] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1816] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1815] = 42'b100000000000000000000010010000000000000000;
    n1466[1814] = 42'b100000000000000000000010110010000000000000;
    n1466[1813] = 42'b000000000000000000000000000110000000000000;
    n1466[1812] = 42'b100000000000000000000000000000010000000100;
    n1466[1811] = 42'b000000000000000000000001110000000000000000;
    n1466[1810] = 42'b100000001001010000000000000000010010001100;
    n1466[1809] = 42'b101000000000000000000000000000000000001110;
    n1466[1808] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1807] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1806] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1805] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1804] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1803] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1802] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1801] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1800] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1799] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1798] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1797] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1796] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1795] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1794] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1793] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1792] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1791] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1790] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1789] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1788] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1787] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1786] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1785] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1784] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1783] = 42'b100000000000000000000010010000000000000000;
    n1466[1782] = 42'b000000000000000000000000110000000000000000;
    n1466[1781] = 42'b100000000000000000000000100000000000001100;
    n1466[1780] = 42'b100000000000000000000001010010000000001100;
    n1466[1779] = 42'b000000000000000000000000000000000000000000;
    n1466[1778] = 42'b100000000000000000000000000000010000000100;
    n1466[1777] = 42'b000000000000000000000001110000000000000000;
    n1466[1776] = 42'b100000000101010000000000000000010010001100;
    n1466[1775] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1774] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1773] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1772] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1771] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1770] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1769] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1768] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1767] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1766] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1765] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1764] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1763] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1762] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1761] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1760] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1759] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1758] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1757] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1756] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1755] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1754] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1753] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1752] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1751] = 42'b100000000000000000000010010000000000000000;
    n1466[1750] = 42'b000000000000000000000000000000000000000000;
    n1466[1749] = 42'b100000000000000000000000000000010000001100;
    n1466[1748] = 42'b000000000000000000000001110000000000000000;
    n1466[1747] = 42'b100000000101010000000000000000010010001100;
    n1466[1746] = 42'b101000000000000000000000000000000000001110;
    n1466[1745] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1744] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1743] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1742] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1741] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1740] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1739] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1738] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1737] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1736] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1735] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1734] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1733] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1732] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1731] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1730] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1729] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1728] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1727] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1726] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1725] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1724] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1723] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1722] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1721] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1720] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1719] = 42'b100000000000000000000010000000010000000000;
    n1466[1718] = 42'b000000000000000000000001110000000000000000;
    n1466[1717] = 42'b100000000101010000000000000000010010001100;
    n1466[1716] = 42'b101000000000000000000000000000000000001110;
    n1466[1715] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1714] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1713] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1712] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1711] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1710] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1709] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1708] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1707] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1706] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1705] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1704] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1703] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1702] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1701] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1700] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1699] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1698] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1697] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1696] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1695] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1694] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1693] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1692] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1691] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1690] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1689] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1688] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1687] = 42'b100000000000000000000010010000000000000000;
    n1466[1686] = 42'b100000000000000000000010000010000000000000;
    n1466[1685] = 42'b000000000000000000000000000000000000000000;
    n1466[1684] = 42'b100000000000000000000000000000010000000100;
    n1466[1683] = 42'b000000000000000000000001110000000000000000;
    n1466[1682] = 42'b100000000101010000000000000000010010001100;
    n1466[1681] = 42'b101000000000000000000000000000000000001110;
    n1466[1680] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1679] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1678] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1677] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1676] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1675] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1674] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1673] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1672] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1671] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1670] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1669] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1668] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1667] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1666] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1665] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1664] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1663] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1662] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1661] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1660] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1659] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1658] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1657] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1656] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1655] = 42'b100000000000000000000010010000000000000000;
    n1466[1654] = 42'b000000000000000000000000000000000000000000;
    n1466[1653] = 42'b100000000000000000000000100000000000001100;
    n1466[1652] = 42'b100000000000000000000001100010000000001100;
    n1466[1651] = 42'b000000000000000000000000000110000000000000;
    n1466[1650] = 42'b100000000000000000000000000000010000000100;
    n1466[1649] = 42'b000000000000000000000001110000000000000000;
    n1466[1648] = 42'b100000000101010000000000000000010010001100;
    n1466[1647] = 42'b100000000000000000000010010000000000000000;
    n1466[1646] = 42'b000000000000000000000000000000000000000000;
    n1466[1645] = 42'b100000000000000000000000100000000000001100;
    n1466[1644] = 42'b100000000000000000000001010010000000001100;
    n1466[1643] = 42'b000000000000000000000000000000000000000000;
    n1466[1642] = 42'b100000000000000000000000000000010000000100;
    n1466[1641] = 42'b000000000000000000000001110000000000000000;
    n1466[1640] = 42'b100000000101010000000000000000010010001100;
    n1466[1639] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1638] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1637] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1636] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1635] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1634] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1633] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1632] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1631] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1630] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1629] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1628] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1627] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1626] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1625] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1624] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1623] = 42'b100000000000000000000010010000000000000000;
    n1466[1622] = 42'b000000000000000000000000110000000000000000;
    n1466[1621] = 42'b100000000000000000000000000000010000001100;
    n1466[1620] = 42'b000000000000000000000001110000000000000000;
    n1466[1619] = 42'b100000000101010000000000000000010010001100;
    n1466[1618] = 42'b101000000000000000000000000000000000001110;
    n1466[1617] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1616] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1615] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1614] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1613] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1612] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1611] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1610] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1609] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1608] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1607] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1606] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1605] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1604] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1603] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1602] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1601] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1600] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1599] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1598] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1597] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1596] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1595] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1594] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1593] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1592] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1591] = 42'b100000000000000000000010010000000000000000;
    n1466[1590] = 42'b100000000000000000000011000010000000000000;
    n1466[1589] = 42'b000000000000000000000000000110000000000000;
    n1466[1588] = 42'b100000000000000000000000000000010000000100;
    n1466[1587] = 42'b000000000000000000000001110000000000000000;
    n1466[1586] = 42'b100000000101010000000000000000010010001100;
    n1466[1585] = 42'b101000000000000000000000000000000000001110;
    n1466[1584] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1583] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1582] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1581] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1580] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1579] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1578] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1577] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1576] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1575] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1574] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1573] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1572] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1571] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1570] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1569] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1568] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1567] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1566] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1565] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1564] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1563] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1562] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1561] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1560] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1559] = 42'b100000000000000000000010010000000000000000;
    n1466[1558] = 42'b100000000000000000000010110010000000000000;
    n1466[1557] = 42'b000000000000000000000000000110000000000000;
    n1466[1556] = 42'b100000000000000000000000000000010000000100;
    n1466[1555] = 42'b000000000000000000000001110000000000000000;
    n1466[1554] = 42'b100000000101010000000000000000010010001100;
    n1466[1553] = 42'b101000000000000000000000000000000000001110;
    n1466[1552] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1551] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1550] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1549] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1548] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1547] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1546] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1545] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1544] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1543] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1542] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1541] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1540] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1539] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1538] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1537] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1536] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1535] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1534] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1533] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1532] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1531] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1530] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1529] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1528] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1527] = 42'b100000000000000000000010010000000000000000;
    n1466[1526] = 42'b000000000000000000000000110000000000000000;
    n1466[1525] = 42'b100000000000000000000000100000000000001100;
    n1466[1524] = 42'b100000000000000000000001010010000000001100;
    n1466[1523] = 42'b000000000000000000000000000000000000000000;
    n1466[1522] = 42'b100000000000000000000000000000010000000100;
    n1466[1521] = 42'b000000000000000000000001110000000000000000;
    n1466[1520] = 42'b100000001101010000000000000000010010001100;
    n1466[1519] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1518] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1517] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1516] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1515] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1514] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1513] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1512] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1511] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1510] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1509] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1508] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1507] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1506] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1505] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1504] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1503] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1502] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1501] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1500] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1499] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1498] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1497] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1496] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1495] = 42'b100000000000000000000010010000000000000000;
    n1466[1494] = 42'b000000000000000000000000000000000000000000;
    n1466[1493] = 42'b100000000000000000000000000000010000001100;
    n1466[1492] = 42'b000000000000000000000001110000000000000000;
    n1466[1491] = 42'b100000001101010000000000000000010010001100;
    n1466[1490] = 42'b101000000000000000000000000000000000001110;
    n1466[1489] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1488] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1487] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1486] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1485] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1484] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1483] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1482] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1481] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1480] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1479] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1478] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1477] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1476] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1475] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1474] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1473] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1472] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1471] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1470] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1469] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1468] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1467] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1466] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1465] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1464] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1463] = 42'b100000000000000000000010000000010000000000;
    n1466[1462] = 42'b000000000000000000000001110000000000000000;
    n1466[1461] = 42'b100000001101010000000000000000010010001100;
    n1466[1460] = 42'b101000000000000000000000000000000000001110;
    n1466[1459] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1458] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1457] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1456] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1455] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1454] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1453] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1452] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1451] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1450] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1449] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1448] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1447] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1446] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1445] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1444] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1443] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1442] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1441] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1440] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1439] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1438] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1437] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1436] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1435] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1434] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1433] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1432] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1431] = 42'b100000000000000000000010010000000000000000;
    n1466[1430] = 42'b100000000000000000000010000010000000000000;
    n1466[1429] = 42'b000000000000000000000000000000000000000000;
    n1466[1428] = 42'b100000000000000000000000000000010000000100;
    n1466[1427] = 42'b000000000000000000000001110000000000000000;
    n1466[1426] = 42'b100000001101010000000000000000010010001100;
    n1466[1425] = 42'b101000000000000000000000000000000000001110;
    n1466[1424] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1423] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1422] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1421] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1420] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1419] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1418] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1417] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1416] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1415] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1414] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1413] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1412] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1411] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1410] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1409] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1408] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1407] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1406] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1405] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1404] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1403] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1402] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1401] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1400] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1399] = 42'b100000000000000000000010010000000000000000;
    n1466[1398] = 42'b000000000000000000000000000000000000000000;
    n1466[1397] = 42'b100000000000000000000000100000000000001100;
    n1466[1396] = 42'b100000000000000000000001100010000000001100;
    n1466[1395] = 42'b000000000000000000000000000110000000000000;
    n1466[1394] = 42'b100000000000000000000000000000010000000100;
    n1466[1393] = 42'b000000000000000000000001110000000000000000;
    n1466[1392] = 42'b100000001101010000000000000000010010001100;
    n1466[1391] = 42'b100000000000000000000010010000000000000000;
    n1466[1390] = 42'b000000000000000000000000000000000000000000;
    n1466[1389] = 42'b100000000000000000000000100000000000001100;
    n1466[1388] = 42'b100000000000000000000001010010000000001100;
    n1466[1387] = 42'b000000000000000000000000000000000000000000;
    n1466[1386] = 42'b100000000000000000000000000000010000000100;
    n1466[1385] = 42'b000000000000000000000001110000000000000000;
    n1466[1384] = 42'b100000001101010000000000000000010010001100;
    n1466[1383] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1382] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1381] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1380] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1379] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1378] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1377] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1376] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1375] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1374] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1373] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1372] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1371] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1370] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1369] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1368] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1367] = 42'b100000000000000000000010010000000000000000;
    n1466[1366] = 42'b000000000000000000000000110000000000000000;
    n1466[1365] = 42'b100000000000000000000000000000010000001100;
    n1466[1364] = 42'b000000000000000000000001110000000000000000;
    n1466[1363] = 42'b100000001101010000000000000000010010001100;
    n1466[1362] = 42'b101000000000000000000000000000000000001110;
    n1466[1361] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1360] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1359] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1358] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1357] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1356] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1355] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1354] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1353] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1352] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1351] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1350] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1349] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1348] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1347] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1346] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1345] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1344] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1343] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1342] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1341] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1340] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1339] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1338] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1337] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1336] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1335] = 42'b100000000000000000000010010000000000000000;
    n1466[1334] = 42'b100000000000000000000011000010000000000000;
    n1466[1333] = 42'b000000000000000000000000000110000000000000;
    n1466[1332] = 42'b100000000000000000000000000000010000000100;
    n1466[1331] = 42'b000000000000000000000001110000000000000000;
    n1466[1330] = 42'b100000001101010000000000000000010010001100;
    n1466[1329] = 42'b101000000000000000000000000000000000001110;
    n1466[1328] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1327] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1326] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1325] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1324] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1323] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1322] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1321] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1320] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1319] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1318] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1317] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1316] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1315] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1314] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1313] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1312] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1311] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1310] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1309] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1308] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1307] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1306] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1305] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1304] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1303] = 42'b100000000000000000000010010000000000000000;
    n1466[1302] = 42'b100000000000000000000010110010000000000000;
    n1466[1301] = 42'b000000000000000000000000000110000000000000;
    n1466[1300] = 42'b100000000000000000000000000000010000000100;
    n1466[1299] = 42'b000000000000000000000001110000000000000000;
    n1466[1298] = 42'b100000001101010000000000000000010010001100;
    n1466[1297] = 42'b101000000000000000000000000000000000001110;
    n1466[1296] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1295] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1294] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1293] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1292] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1291] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1290] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1289] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1288] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1287] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1286] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1285] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1284] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1283] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1282] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1281] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1280] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1279] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1278] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1277] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1276] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1275] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1274] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1273] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1272] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1271] = 42'b100000000000000000000010010000000000000000;
    n1466[1270] = 42'b000000000000000000000000110000000000000000;
    n1466[1269] = 42'b100000000000000000000000100000000000001100;
    n1466[1268] = 42'b100000000000000000000001010010000000001100;
    n1466[1267] = 42'b000000000000000000000000000000000000000000;
    n1466[1266] = 42'b100000000000000000000000000000010000000100;
    n1466[1265] = 42'b000000000000000000000001110000000000000000;
    n1466[1264] = 42'b100000010001010000000000000000011010001100;
    n1466[1263] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1262] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1261] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1260] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1259] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1258] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1257] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1256] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1255] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1254] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1253] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1252] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1251] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1250] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1249] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1248] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1247] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1246] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1245] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1244] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1243] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1242] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1241] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1240] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1239] = 42'b100000000000000000000010010000000000000000;
    n1466[1238] = 42'b000000000000000000000000000000000000000000;
    n1466[1237] = 42'b100000000000000000000000000000010000001100;
    n1466[1236] = 42'b000000000000000000000001110000000000000000;
    n1466[1235] = 42'b100000010001010000000000000000011010001100;
    n1466[1234] = 42'b101000000000000000000000000000000000001101;
    n1466[1233] = 42'b000000000000000000000000000000000000000010;
    n1466[1232] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1231] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1230] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1229] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1228] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1227] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1226] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1225] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1224] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1223] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1222] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1221] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1220] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1219] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1218] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1217] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1216] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1215] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1214] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1213] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1212] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1211] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1210] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1209] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1208] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1207] = 42'b100000000000000000000010000000010000000000;
    n1466[1206] = 42'b000000000000000000000001110000000000000000;
    n1466[1205] = 42'b100000010001010000000000000000011010001100;
    n1466[1204] = 42'b101000000000000000000000000000000000001101;
    n1466[1203] = 42'b000000000000000000000000000000000000000010;
    n1466[1202] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1201] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1200] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1199] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1198] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1197] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1196] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1195] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1194] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1193] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1192] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1191] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1190] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1189] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1188] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1187] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1186] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1185] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1184] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1183] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1182] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1181] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1180] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1179] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1178] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1177] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1176] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1175] = 42'b100000000000000000000010010000000000000000;
    n1466[1174] = 42'b100000000000000000000010000010000000000000;
    n1466[1173] = 42'b000000000000000000000000000000000000000000;
    n1466[1172] = 42'b100000000000000000000000000000010000000100;
    n1466[1171] = 42'b000000000000000000000001110000000000000000;
    n1466[1170] = 42'b100000010001010000000000000000011010001100;
    n1466[1169] = 42'b101000000000000000000000000000000000001101;
    n1466[1168] = 42'b000000000000000000000000000000000000000010;
    n1466[1167] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1166] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1165] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1164] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1163] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1162] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1161] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1160] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1159] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1158] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1157] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1156] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1155] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1154] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1153] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1152] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1151] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1150] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1149] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1148] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1147] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1146] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1145] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1144] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1143] = 42'b100000000000000000000010010000000000000000;
    n1466[1142] = 42'b000000000000000000000000000000000000000000;
    n1466[1141] = 42'b100000000000000000000000100000000000001100;
    n1466[1140] = 42'b100000000000000000000001100010000000001100;
    n1466[1139] = 42'b000000000000000000000000000110000000000000;
    n1466[1138] = 42'b100000000000000000000000000000010000000100;
    n1466[1137] = 42'b000000000000000000000001110000000000000000;
    n1466[1136] = 42'b100000010001010000000000000000011010001100;
    n1466[1135] = 42'b100000000000000000000010010000000000000000;
    n1466[1134] = 42'b000000000000000000000000000000000000000000;
    n1466[1133] = 42'b100000000000000000000000100000000000001100;
    n1466[1132] = 42'b100000000000000000000001010010000000001100;
    n1466[1131] = 42'b000000000000000000000000000000000000000000;
    n1466[1130] = 42'b100000000000000000000000000000010000000100;
    n1466[1129] = 42'b000000000000000000000001110000000000000000;
    n1466[1128] = 42'b100000010001010000000000000000011010001100;
    n1466[1127] = 42'b100000000000000010000010000000000000000000;
    n1466[1126] = 42'b100000000000000000000010000000000001100000;
    n1466[1125] = 42'b000000000000000000000000000000000000000000;
    n1466[1124] = 42'b000000000000000000000000000000000000000000;
    n1466[1123] = 42'b000000011000010000000000000000000000000000;
    n1466[1122] = 42'b000001000010100000000000000000000000000000;
    n1466[1121] = 42'b100000011100100100000000000001000000011000;
    n1466[1120] = 42'b000001000110000000000000000000000000100000;
    n1466[1119] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1118] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1117] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1116] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1115] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1114] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1113] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1112] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1111] = 42'b100000000000000000000010010000000000000000;
    n1466[1110] = 42'b000000000000000000000000110000000000000000;
    n1466[1109] = 42'b100000000000000000000000000000010000001100;
    n1466[1108] = 42'b000000000000000000000001110000000000000000;
    n1466[1107] = 42'b100000010001010000000000000000011010001100;
    n1466[1106] = 42'b101000000000000000000000000000000000001101;
    n1466[1105] = 42'b000000000000000000000000000000000000000010;
    n1466[1104] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1103] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1102] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1101] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1100] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1099] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1098] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1097] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1096] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1095] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1094] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1093] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1092] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1091] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1090] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1089] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1088] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1087] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1086] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1085] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1084] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1083] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1082] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1081] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1080] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1079] = 42'b100000000000000000000010010000000000000000;
    n1466[1078] = 42'b100000000000000000000011000010000000000000;
    n1466[1077] = 42'b000000000000000000000000000110000000000000;
    n1466[1076] = 42'b100000000000000000000000000000010000000100;
    n1466[1075] = 42'b000000000000000000000001110000000000000000;
    n1466[1074] = 42'b100000010001010000000000000000011010001100;
    n1466[1073] = 42'b101000000000000000000000000000000000001101;
    n1466[1072] = 42'b000000000000000000000000000000000000000010;
    n1466[1071] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1070] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1069] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1068] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1067] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1066] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1065] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1064] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1063] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1062] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1061] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1060] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1059] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1058] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1057] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1056] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1055] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1054] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1053] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1052] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1051] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1050] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1049] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1048] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1047] = 42'b100000000000000000000010010000000000000000;
    n1466[1046] = 42'b100000000000000000000010110010000000000000;
    n1466[1045] = 42'b000000000000000000000000000110000000000000;
    n1466[1044] = 42'b100000000000000000000000000000010000000100;
    n1466[1043] = 42'b000000000000000000000001110000000000000000;
    n1466[1042] = 42'b100000010001010000000000000000011010001100;
    n1466[1041] = 42'b101000000000000000000000000000000000001101;
    n1466[1040] = 42'b000000000000000000000000000000000000000010;
    n1466[1039] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1038] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1037] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1036] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1035] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1034] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1033] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1032] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1031] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1030] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1029] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1028] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1027] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1026] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1025] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1024] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1023] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1022] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1021] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1020] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1019] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1018] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1017] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1016] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1015] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1014] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1013] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1012] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1011] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1010] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1009] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1008] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1007] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1006] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1005] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1004] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1003] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1002] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1001] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1000] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[999] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[998] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[997] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[996] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[995] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[994] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[993] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[992] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[991] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[990] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[989] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[988] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[987] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[986] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[985] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[984] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[983] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[982] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[981] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[980] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[979] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[978] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[977] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[976] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[975] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[974] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[973] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[972] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[971] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[970] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[969] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[968] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[967] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[966] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[965] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[964] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[963] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[962] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[961] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[960] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[959] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[958] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[957] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[956] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[955] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[954] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[953] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[952] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[951] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[950] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[949] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[948] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[947] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[946] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[945] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[944] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[943] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[942] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[941] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[940] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[939] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[938] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[937] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[936] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[935] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[934] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[933] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[932] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[931] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[930] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[929] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[928] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[927] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[926] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[925] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[924] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[923] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[922] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[921] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[920] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[919] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[918] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[917] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[916] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[915] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[914] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[913] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[912] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[911] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[910] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[909] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[908] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[907] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[906] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[905] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[904] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[903] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[902] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[901] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[900] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[899] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[898] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[897] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[896] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[895] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[894] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[893] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[892] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[891] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[890] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[889] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[888] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[887] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[886] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[885] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[884] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[883] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[882] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[881] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[880] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[879] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[878] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[877] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[876] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[875] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[874] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[873] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[872] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[871] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[870] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[869] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[868] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[867] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[866] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[865] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[864] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[863] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[862] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[861] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[860] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[859] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[858] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[857] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[856] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[855] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[854] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[853] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[852] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[851] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[850] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[849] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[848] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[847] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[846] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[845] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[844] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[843] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[842] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[841] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[840] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[839] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[838] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[837] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[836] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[835] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[834] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[833] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[832] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[831] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[830] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[829] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[828] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[827] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[826] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[825] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[824] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[823] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[822] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[821] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[820] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[819] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[818] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[817] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[816] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[815] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[814] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[813] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[812] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[811] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[810] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[809] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[808] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[807] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[806] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[805] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[804] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[803] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[802] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[801] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[800] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[799] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[798] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[797] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[796] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[795] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[794] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[793] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[792] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[791] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[790] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[789] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[788] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[787] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[786] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[785] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[784] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[783] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[782] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[781] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[780] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[779] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[778] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[777] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[776] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[775] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[774] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[773] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[772] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[771] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[770] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[769] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[768] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[767] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[766] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[765] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[764] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[763] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[762] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[761] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[760] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[759] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[758] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[757] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[756] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[755] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[754] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[753] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[752] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[751] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[750] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[749] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[748] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[747] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[746] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[745] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[744] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[743] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[742] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[741] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[740] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[739] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[738] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[737] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[736] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[735] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[734] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[733] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[732] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[731] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[730] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[729] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[728] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[727] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[726] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[725] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[724] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[723] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[722] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[721] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[720] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[719] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[718] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[717] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[716] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[715] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[714] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[713] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[712] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[711] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[710] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[709] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[708] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[707] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[706] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[705] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[704] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[703] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[702] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[701] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[700] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[699] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[698] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[697] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[696] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[695] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[694] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[693] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[692] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[691] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[690] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[689] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[688] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[687] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[686] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[685] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[684] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[683] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[682] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[681] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[680] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[679] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[678] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[677] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[676] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[675] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[674] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[673] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[672] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[671] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[670] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[669] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[668] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[667] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[666] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[665] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[664] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[663] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[662] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[661] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[660] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[659] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[658] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[657] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[656] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[655] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[654] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[653] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[652] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[651] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[650] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[649] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[648] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[647] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[646] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[645] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[644] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[643] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[642] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[641] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[640] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[639] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[638] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[637] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[636] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[635] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[634] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[633] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[632] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[631] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[630] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[629] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[628] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[627] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[626] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[625] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[624] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[623] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[622] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[621] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[620] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[619] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[618] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[617] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[616] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[615] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[614] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[613] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[612] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[611] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[610] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[609] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[608] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[607] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[606] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[605] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[604] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[603] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[602] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[601] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[600] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[599] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[598] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[597] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[596] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[595] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[594] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[593] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[592] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[591] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[590] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[589] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[588] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[587] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[586] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[585] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[584] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[583] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[582] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[581] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[580] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[579] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[578] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[577] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[576] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[575] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[574] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[573] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[572] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[571] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[570] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[569] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[568] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[567] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[566] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[565] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[564] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[563] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[562] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[561] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[560] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[559] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[558] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[557] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[556] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[555] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[554] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[553] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[552] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[551] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[550] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[549] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[548] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[547] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[546] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[545] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[544] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[543] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[542] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[541] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[540] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[539] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[538] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[537] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[536] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[535] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[534] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[533] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[532] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[531] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[530] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[529] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[528] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[527] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[526] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[525] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[524] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[523] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[522] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[521] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[520] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[519] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[518] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[517] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[516] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[515] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[514] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[513] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[512] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[511] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[510] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[509] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[508] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[507] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[506] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[505] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[504] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[503] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[502] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[501] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[500] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[499] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[498] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[497] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[496] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[495] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[494] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[493] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[492] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[491] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[490] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[489] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[488] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[487] = 42'b100000000000000010000010000000000000000000;
    n1466[486] = 42'b100000000000000000000010000000000001100000;
    n1466[485] = 42'b000000000000000000000000000000000000000000;
    n1466[484] = 42'b000000000000000000000000000000000000000000;
    n1466[483] = 42'b000000011000010000000000000000000000000000;
    n1466[482] = 42'b000001000010100000000000000000000000000000;
    n1466[481] = 42'b100000011000100100000000000001000000011000;
    n1466[480] = 42'b000001000010000000000000000000000000100000;
    n1466[479] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[478] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[477] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[476] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[475] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[474] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[473] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[472] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[471] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[470] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[469] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[468] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[467] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[466] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[465] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[464] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[463] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[462] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[461] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[460] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[459] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[458] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[457] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[456] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[455] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[454] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[453] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[452] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[451] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[450] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[449] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[448] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[447] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[446] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[445] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[444] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[443] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[442] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[441] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[440] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[439] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[438] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[437] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[436] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[435] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[434] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[433] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[432] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[431] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[430] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[429] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[428] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[427] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[426] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[425] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[424] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[423] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[422] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[421] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[420] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[419] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[418] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[417] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[416] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[415] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[414] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[413] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[412] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[411] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[410] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[409] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[408] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[407] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[406] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[405] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[404] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[403] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[402] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[401] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[400] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[399] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[398] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[397] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[396] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[395] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[394] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[393] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[392] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[391] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[390] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[389] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[388] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[387] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[386] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[385] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[384] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[383] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[382] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[381] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[380] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[379] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[378] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[377] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[376] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[375] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[374] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[373] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[372] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[371] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[370] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[369] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[368] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[367] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[366] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[365] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[364] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[363] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[362] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[361] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[360] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[359] = 42'b100000000000000010000010000000000000000000;
    n1466[358] = 42'b100000000000000000000010000000000001100000;
    n1466[357] = 42'b000000000000000000000000000000000000000000;
    n1466[356] = 42'b000000000000000000000000000000000000000000;
    n1466[355] = 42'b000000011000010000000000000000000000000000;
    n1466[354] = 42'b000001000010100000000000000000000000000000;
    n1466[353] = 42'b100000011100100100000000000001000000011000;
    n1466[352] = 42'b000001000110000000000000000000000000100000;
    n1466[351] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[350] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[349] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[348] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[347] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[346] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[345] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[344] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[343] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[342] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[341] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[340] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[339] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[338] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[337] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[336] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[335] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[334] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[333] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[332] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[331] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[330] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[329] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[328] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[327] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[326] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[325] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[324] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[323] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[322] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[321] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[320] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[319] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[318] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[317] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[316] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[315] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[314] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[313] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[312] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[311] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[310] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[309] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[308] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[307] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[306] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[305] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[304] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[303] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[302] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[301] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[300] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[299] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[298] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[297] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[296] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[295] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[294] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[293] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[292] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[291] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[290] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[289] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[288] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[287] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[286] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[285] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[284] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[283] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[282] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[281] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[280] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[279] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[278] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[277] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[276] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[275] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[274] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[273] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[272] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[271] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[270] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[269] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[268] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[267] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[266] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[265] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[264] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[263] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[262] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[261] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[260] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[259] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[258] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[257] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[256] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[255] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[254] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[253] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[252] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[251] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[250] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[249] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[248] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[247] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[246] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[245] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[244] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[243] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[242] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[241] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[240] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[239] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[238] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[237] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[236] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[235] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[234] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[233] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[232] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[231] = 42'b100000000000000010000010000000000000000000;
    n1466[230] = 42'b100000000000000000000010000000000001100000;
    n1466[229] = 42'b000000000000000000000000000000000000000000;
    n1466[228] = 42'b000000000000000000000000000000000000000000;
    n1466[227] = 42'b000000011000010000000000000000000000000000;
    n1466[226] = 42'b000001000010100000000000000000000000000000;
    n1466[225] = 42'b100000011100100100000000000001000000011000;
    n1466[224] = 42'b000001000110000000000000000000000000100000;
    n1466[223] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[222] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[221] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[220] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[219] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[218] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[217] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[216] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[215] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[214] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[213] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[212] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[211] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[210] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[209] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[208] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[207] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[206] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[205] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[204] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[203] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[202] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[201] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[200] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[199] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[198] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[197] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[196] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[195] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[194] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[193] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[192] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[191] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[190] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[189] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[188] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[187] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[186] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[185] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[184] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[183] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[182] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[181] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[180] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[179] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[178] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[177] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[176] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[175] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[174] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[173] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[172] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[171] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[170] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[169] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[168] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[167] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[166] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[165] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[164] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[163] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[162] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[161] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[160] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[159] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[158] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[157] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[156] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[155] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[154] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[153] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[152] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[151] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[150] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[149] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[148] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[147] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[146] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[145] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[144] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[143] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[142] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[141] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[140] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[139] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[138] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[137] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[136] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[135] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[134] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[133] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[132] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[131] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[130] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[129] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[128] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[127] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[126] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[125] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[124] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[123] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[122] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[121] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[120] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[119] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[118] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[117] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[116] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[115] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[114] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[113] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[112] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[111] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[110] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[109] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[108] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[107] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[106] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[105] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[104] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[103] = 42'b100000000000000010000010000000000000000000;
    n1466[102] = 42'b100000000000000000000010000000000001100000;
    n1466[101] = 42'b000000000000000000000000000000000000000000;
    n1466[100] = 42'b000000000000000000000000000000000000000000;
    n1466[99] = 42'b000000011000010000000000000000000000000000;
    n1466[98] = 42'b000001000010100000000000000000000000000000;
    n1466[97] = 42'b100000011000100100000000000001000000011000;
    n1466[96] = 42'b000001000010000000000000000000000000100000;
    n1466[95] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[94] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[93] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[92] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[91] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[90] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[89] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[88] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[87] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[86] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[85] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[84] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[83] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[82] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[81] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[80] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[79] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[78] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[77] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[76] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[75] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[74] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[73] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[72] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[71] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[70] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[69] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[68] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[67] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[66] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[65] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[64] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[63] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[62] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[61] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[60] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[59] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[58] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[57] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[56] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[55] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[54] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[53] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[52] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[51] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[50] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[49] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[48] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[47] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[46] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[45] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[44] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[43] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[42] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[41] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[40] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[39] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[38] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[37] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[36] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[35] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[34] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[33] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[32] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[31] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[30] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[29] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[28] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[27] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[26] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[25] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[24] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[23] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[22] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[21] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[20] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[19] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[18] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[17] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[16] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[15] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[14] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[13] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[12] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[11] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[10] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[9] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[8] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[7] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[6] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[5] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[4] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[3] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[2] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[1] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1466[0] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    end
  assign n1467_data = n1466[n1414_o];
  /* HUC6280_MC.vhd:6986:54  */
  /* HUC6280_MC.vhd:6986:53  */
  reg [41:0] n1468[2047:0] ; // memory
  initial begin
    n1468[2047] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2046] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2045] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2044] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2043] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2042] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2041] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2040] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2039] = 42'b101000000000000000000000000000000000001110;
    n1468[2038] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2037] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2036] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2035] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2034] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2033] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2032] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2031] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2030] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2029] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2028] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2027] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2026] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2025] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2024] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2023] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2022] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2021] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2020] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2019] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2018] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2017] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2016] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2015] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2014] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2013] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2012] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2011] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2010] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2009] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2008] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2007] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2006] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2005] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2004] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2003] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2002] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2001] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2000] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1999] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1998] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1997] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1996] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1995] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1994] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1993] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1992] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1991] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1990] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1989] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1988] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1987] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1986] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1985] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1984] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1983] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1982] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1981] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1980] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1979] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1978] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1977] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1976] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1975] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1974] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1973] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1972] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1971] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1970] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1969] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1968] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1967] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1966] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1965] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1964] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1963] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1962] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1961] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1960] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1959] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1958] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1957] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1956] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1955] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1954] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1953] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1952] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1951] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1950] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1949] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1948] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1947] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1946] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1945] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1944] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1943] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1942] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1941] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1940] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1939] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1938] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1937] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1936] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1935] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1934] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1933] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1932] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1931] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1930] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1929] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1928] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1927] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1926] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1925] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1924] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1923] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1922] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1921] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1920] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1919] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1918] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1917] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1916] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1915] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1914] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1913] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1912] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1911] = 42'b101000000000000000000000000000000000001110;
    n1468[1910] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1909] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1908] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1907] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1906] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1905] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1904] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1903] = 42'b101000000000000000000000000000000000001110;
    n1468[1902] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1901] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1900] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1899] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1898] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1897] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1896] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1895] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1894] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1893] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1892] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1891] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1890] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1889] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1888] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1887] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1886] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1885] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1884] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1883] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1882] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1881] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1880] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1879] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1878] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1877] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1876] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1875] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1874] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1873] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1872] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1871] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1870] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1869] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1868] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1867] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1866] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1865] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1864] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1863] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1862] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1861] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1860] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1859] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1858] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1857] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1856] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1855] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1854] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1853] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1852] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1851] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1850] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1849] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1848] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1847] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1846] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1845] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1844] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1843] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1842] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1841] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1840] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1839] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1838] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1837] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1836] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1835] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1834] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1833] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1832] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1831] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1830] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1829] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1828] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1827] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1826] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1825] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1824] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1823] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1822] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1821] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1820] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1819] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1818] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1817] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1816] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1815] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1814] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1813] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1812] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1811] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1810] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1809] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1808] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1807] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1806] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1805] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1804] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1803] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1802] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1801] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1800] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1799] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1798] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1797] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1796] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1795] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1794] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1793] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1792] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1791] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1790] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1789] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1788] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1787] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1786] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1785] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1784] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1783] = 42'b101000000000000000000000000000000000001110;
    n1468[1782] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1781] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1780] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1779] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1778] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1777] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1776] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1775] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1774] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1773] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1772] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1771] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1770] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1769] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1768] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1767] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1766] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1765] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1764] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1763] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1762] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1761] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1760] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1759] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1758] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1757] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1756] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1755] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1754] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1753] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1752] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1751] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1750] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1749] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1748] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1747] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1746] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1745] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1744] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1743] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1742] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1741] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1740] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1739] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1738] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1737] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1736] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1735] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1734] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1733] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1732] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1731] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1730] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1729] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1728] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1727] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1726] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1725] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1724] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1723] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1722] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1721] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1720] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1719] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1718] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1717] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1716] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1715] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1714] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1713] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1712] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1711] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1710] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1709] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1708] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1707] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1706] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1705] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1704] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1703] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1702] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1701] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1700] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1699] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1698] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1697] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1696] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1695] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1694] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1693] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1692] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1691] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1690] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1689] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1688] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1687] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1686] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1685] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1684] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1683] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1682] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1681] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1680] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1679] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1678] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1677] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1676] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1675] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1674] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1673] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1672] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1671] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1670] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1669] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1668] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1667] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1666] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1665] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1664] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1663] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1662] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1661] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1660] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1659] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1658] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1657] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1656] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1655] = 42'b101000000000000000000000000000000000001110;
    n1468[1654] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1653] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1652] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1651] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1650] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1649] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1648] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1647] = 42'b101000000000000000000000000000000000001110;
    n1468[1646] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1645] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1644] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1643] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1642] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1641] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1640] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1639] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1638] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1637] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1636] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1635] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1634] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1633] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1632] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1631] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1630] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1629] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1628] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1627] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1626] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1625] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1624] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1623] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1622] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1621] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1620] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1619] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1618] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1617] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1616] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1615] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1614] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1613] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1612] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1611] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1610] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1609] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1608] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1607] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1606] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1605] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1604] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1603] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1602] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1601] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1600] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1599] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1598] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1597] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1596] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1595] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1594] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1593] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1592] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1591] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1590] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1589] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1588] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1587] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1586] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1585] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1584] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1583] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1582] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1581] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1580] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1579] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1578] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1577] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1576] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1575] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1574] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1573] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1572] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1571] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1570] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1569] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1568] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1567] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1566] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1565] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1564] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1563] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1562] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1561] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1560] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1559] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1558] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1557] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1556] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1555] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1554] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1553] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1552] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1551] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1550] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1549] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1548] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1547] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1546] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1545] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1544] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1543] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1542] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1541] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1540] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1539] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1538] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1537] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1536] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1535] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1534] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1533] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1532] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1531] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1530] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1529] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1528] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1527] = 42'b101000000000000000000000000000000000001110;
    n1468[1526] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1525] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1524] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1523] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1522] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1521] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1520] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1519] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1518] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1517] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1516] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1515] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1514] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1513] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1512] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1511] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1510] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1509] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1508] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1507] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1506] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1505] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1504] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1503] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1502] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1501] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1500] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1499] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1498] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1497] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1496] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1495] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1494] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1493] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1492] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1491] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1490] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1489] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1488] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1487] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1486] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1485] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1484] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1483] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1482] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1481] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1480] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1479] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1478] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1477] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1476] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1475] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1474] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1473] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1472] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1471] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1470] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1469] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1468] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1467] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1466] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1465] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1464] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1463] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1462] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1461] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1460] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1459] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1458] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1457] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1456] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1455] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1454] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1453] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1452] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1451] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1450] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1449] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1448] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1447] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1446] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1445] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1444] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1443] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1442] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1441] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1440] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1439] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1438] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1437] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1436] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1435] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1434] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1433] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1432] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1431] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1430] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1429] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1428] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1427] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1426] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1425] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1424] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1423] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1422] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1421] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1420] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1419] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1418] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1417] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1416] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1415] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1414] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1413] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1412] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1411] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1410] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1409] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1408] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1407] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1406] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1405] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1404] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1403] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1402] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1401] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1400] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1399] = 42'b101000000000000000000000000000000000001110;
    n1468[1398] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1397] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1396] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1395] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1394] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1393] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1392] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1391] = 42'b101000000000000000000000000000000000001110;
    n1468[1390] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1389] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1388] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1387] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1386] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1385] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1384] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1383] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1382] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1381] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1380] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1379] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1378] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1377] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1376] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1375] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1374] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1373] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1372] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1371] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1370] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1369] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1368] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1367] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1366] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1365] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1364] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1363] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1362] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1361] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1360] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1359] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1358] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1357] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1356] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1355] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1354] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1353] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1352] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1351] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1350] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1349] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1348] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1347] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1346] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1345] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1344] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1343] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1342] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1341] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1340] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1339] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1338] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1337] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1336] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1335] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1334] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1333] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1332] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1331] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1330] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1329] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1328] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1327] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1326] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1325] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1324] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1323] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1322] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1321] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1320] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1319] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1318] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1317] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1316] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1315] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1314] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1313] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1312] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1311] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1310] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1309] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1308] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1307] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1306] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1305] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1304] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1303] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1302] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1301] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1300] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1299] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1298] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1297] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1296] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1295] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1294] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1293] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1292] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1291] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1290] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1289] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1288] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1287] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1286] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1285] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1284] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1283] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1282] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1281] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1280] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1279] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1278] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1277] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1276] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1275] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1274] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1273] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1272] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1271] = 42'b101000000000000000000000000000000000001101;
    n1468[1270] = 42'b000000000000000000000000000000000000000010;
    n1468[1269] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1268] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1267] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1266] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1265] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1264] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1263] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1262] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1261] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1260] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1259] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1258] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1257] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1256] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1255] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1254] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1253] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1252] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1251] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1250] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1249] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1248] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1247] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1246] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1245] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1244] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1243] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1242] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1241] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1240] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1239] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1238] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1237] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1236] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1235] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1234] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1233] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1232] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1231] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1230] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1229] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1228] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1227] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1226] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1225] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1224] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1223] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1222] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1221] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1220] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1219] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1218] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1217] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1216] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1215] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1214] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1213] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1212] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1211] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1210] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1209] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1208] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1207] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1206] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1205] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1204] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1203] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1202] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1201] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1200] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1199] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1198] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1197] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1196] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1195] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1194] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1193] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1192] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1191] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1190] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1189] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1188] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1187] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1186] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1185] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1184] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1183] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1182] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1181] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1180] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1179] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1178] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1177] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1176] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1175] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1174] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1173] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1172] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1171] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1170] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1169] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1168] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1167] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1166] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1165] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1164] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1163] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1162] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1161] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1160] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1159] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1158] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1157] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1156] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1155] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1154] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1153] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1152] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1151] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1150] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1149] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1148] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1147] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1146] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1145] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1144] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1143] = 42'b101000000000000000000000000000000000001101;
    n1468[1142] = 42'b000000000000000000000000000000000000000010;
    n1468[1141] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1140] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1139] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1138] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1137] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1136] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1135] = 42'b101000000000000000000000000000000000001101;
    n1468[1134] = 42'b100000000000000000000000000000000000000010;
    n1468[1133] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1132] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1131] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1130] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1129] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1128] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1127] = 42'b101000011100111000000000000000000000011100;
    n1468[1126] = 42'b000001000110010000000000000000000001000000;
    n1468[1125] = 42'b000000011000010010000000000000000000000000;
    n1468[1124] = 42'b000001000010100000000000000000000001100011;
    n1468[1123] = 42'b100000000000000100100000000000000000001000;
    n1468[1122] = 42'b100000000000000010100000000000000000001000;
    n1468[1121] = 42'b100000000000001000000000000000000000001010;
    n1468[1120] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1119] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1118] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1117] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1116] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1115] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1114] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1113] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1112] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1111] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1110] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1109] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1108] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1107] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1106] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1105] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1104] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1103] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1102] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1101] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1100] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1099] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1098] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1097] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1096] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1095] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1094] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1093] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1092] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1091] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1090] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1089] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1088] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1087] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1086] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1085] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1084] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1083] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1082] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1081] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1080] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1079] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1078] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1077] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1076] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1075] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1074] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1073] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1072] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1071] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1070] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1069] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1068] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1067] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1066] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1065] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1064] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1063] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1062] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1061] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1060] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1059] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1058] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1057] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1056] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1055] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1054] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1053] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1052] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1051] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1050] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1049] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1048] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1047] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1046] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1045] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1044] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1043] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1042] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1041] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1040] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1039] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1038] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1037] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1036] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1035] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1034] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1033] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1032] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1031] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1030] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1029] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1028] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1027] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1026] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1025] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1024] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1023] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1022] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1021] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1020] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1019] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1018] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1017] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1016] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1015] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1014] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1013] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1012] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1011] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1010] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1009] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1008] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1007] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1006] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1005] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1004] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1003] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1002] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1001] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1000] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[999] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[998] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[997] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[996] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[995] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[994] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[993] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[992] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[991] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[990] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[989] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[988] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[987] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[986] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[985] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[984] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[983] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[982] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[981] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[980] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[979] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[978] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[977] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[976] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[975] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[974] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[973] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[972] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[971] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[970] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[969] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[968] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[967] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[966] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[965] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[964] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[963] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[962] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[961] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[960] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[959] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[958] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[957] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[956] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[955] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[954] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[953] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[952] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[951] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[950] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[949] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[948] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[947] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[946] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[945] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[944] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[943] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[942] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[941] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[940] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[939] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[938] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[937] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[936] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[935] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[934] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[933] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[932] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[931] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[930] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[929] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[928] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[927] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[926] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[925] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[924] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[923] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[922] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[921] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[920] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[919] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[918] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[917] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[916] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[915] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[914] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[913] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[912] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[911] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[910] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[909] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[908] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[907] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[906] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[905] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[904] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[903] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[902] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[901] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[900] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[899] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[898] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[897] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[896] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[895] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[894] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[893] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[892] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[891] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[890] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[889] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[888] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[887] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[886] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[885] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[884] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[883] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[882] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[881] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[880] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[879] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[878] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[877] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[876] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[875] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[874] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[873] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[872] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[871] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[870] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[869] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[868] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[867] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[866] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[865] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[864] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[863] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[862] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[861] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[860] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[859] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[858] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[857] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[856] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[855] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[854] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[853] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[852] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[851] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[850] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[849] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[848] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[847] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[846] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[845] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[844] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[843] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[842] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[841] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[840] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[839] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[838] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[837] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[836] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[835] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[834] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[833] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[832] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[831] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[830] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[829] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[828] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[827] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[826] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[825] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[824] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[823] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[822] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[821] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[820] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[819] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[818] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[817] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[816] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[815] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[814] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[813] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[812] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[811] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[810] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[809] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[808] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[807] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[806] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[805] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[804] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[803] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[802] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[801] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[800] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[799] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[798] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[797] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[796] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[795] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[794] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[793] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[792] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[791] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[790] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[789] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[788] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[787] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[786] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[785] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[784] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[783] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[782] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[781] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[780] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[779] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[778] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[777] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[776] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[775] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[774] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[773] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[772] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[771] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[770] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[769] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[768] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[767] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[766] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[765] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[764] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[763] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[762] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[761] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[760] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[759] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[758] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[757] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[756] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[755] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[754] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[753] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[752] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[751] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[750] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[749] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[748] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[747] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[746] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[745] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[744] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[743] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[742] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[741] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[740] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[739] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[738] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[737] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[736] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[735] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[734] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[733] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[732] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[731] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[730] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[729] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[728] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[727] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[726] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[725] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[724] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[723] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[722] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[721] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[720] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[719] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[718] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[717] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[716] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[715] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[714] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[713] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[712] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[711] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[710] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[709] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[708] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[707] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[706] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[705] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[704] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[703] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[702] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[701] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[700] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[699] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[698] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[697] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[696] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[695] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[694] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[693] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[692] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[691] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[690] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[689] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[688] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[687] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[686] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[685] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[684] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[683] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[682] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[681] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[680] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[679] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[678] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[677] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[676] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[675] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[674] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[673] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[672] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[671] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[670] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[669] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[668] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[667] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[666] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[665] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[664] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[663] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[662] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[661] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[660] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[659] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[658] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[657] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[656] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[655] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[654] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[653] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[652] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[651] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[650] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[649] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[648] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[647] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[646] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[645] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[644] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[643] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[642] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[641] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[640] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[639] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[638] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[637] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[636] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[635] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[634] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[633] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[632] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[631] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[630] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[629] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[628] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[627] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[626] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[625] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[624] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[623] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[622] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[621] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[620] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[619] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[618] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[617] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[616] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[615] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[614] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[613] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[612] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[611] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[610] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[609] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[608] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[607] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[606] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[605] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[604] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[603] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[602] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[601] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[600] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[599] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[598] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[597] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[596] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[595] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[594] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[593] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[592] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[591] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[590] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[589] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[588] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[587] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[586] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[585] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[584] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[583] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[582] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[581] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[580] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[579] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[578] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[577] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[576] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[575] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[574] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[573] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[572] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[571] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[570] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[569] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[568] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[567] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[566] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[565] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[564] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[563] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[562] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[561] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[560] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[559] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[558] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[557] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[556] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[555] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[554] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[553] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[552] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[551] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[550] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[549] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[548] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[547] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[546] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[545] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[544] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[543] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[542] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[541] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[540] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[539] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[538] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[537] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[536] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[535] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[534] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[533] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[532] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[531] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[530] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[529] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[528] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[527] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[526] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[525] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[524] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[523] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[522] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[521] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[520] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[519] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[518] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[517] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[516] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[515] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[514] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[513] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[512] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[511] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[510] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[509] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[508] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[507] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[506] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[505] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[504] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[503] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[502] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[501] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[500] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[499] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[498] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[497] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[496] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[495] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[494] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[493] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[492] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[491] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[490] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[489] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[488] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[487] = 42'b101000011000111000000000000000000000011100;
    n1468[486] = 42'b000001000010010000000000000000000001000000;
    n1468[485] = 42'b000000011000010010000000000000000000000000;
    n1468[484] = 42'b000001000010100000000000000000000001100011;
    n1468[483] = 42'b100000000000000100100000000000000000001000;
    n1468[482] = 42'b100000000000000010100000000000000000001000;
    n1468[481] = 42'b100000000000001000000000000000000000001010;
    n1468[480] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[479] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[478] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[477] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[476] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[475] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[474] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[473] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[472] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[471] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[470] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[469] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[468] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[467] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[466] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[465] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[464] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[463] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[462] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[461] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[460] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[459] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[458] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[457] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[456] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[455] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[454] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[453] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[452] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[451] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[450] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[449] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[448] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[447] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[446] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[445] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[444] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[443] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[442] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[441] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[440] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[439] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[438] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[437] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[436] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[435] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[434] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[433] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[432] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[431] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[430] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[429] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[428] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[427] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[426] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[425] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[424] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[423] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[422] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[421] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[420] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[419] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[418] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[417] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[416] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[415] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[414] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[413] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[412] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[411] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[410] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[409] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[408] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[407] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[406] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[405] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[404] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[403] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[402] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[401] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[400] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[399] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[398] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[397] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[396] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[395] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[394] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[393] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[392] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[391] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[390] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[389] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[388] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[387] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[386] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[385] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[384] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[383] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[382] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[381] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[380] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[379] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[378] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[377] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[376] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[375] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[374] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[373] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[372] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[371] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[370] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[369] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[368] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[367] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[366] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[365] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[364] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[363] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[362] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[361] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[360] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[359] = 42'b101000000000000000000000000000000000011100;
    n1468[358] = 42'b000000000000000000000000000000000000000000;
    n1468[357] = 42'b000000011000010010000000000000000000000000;
    n1468[356] = 42'b000001000010100000000000000000000001100011;
    n1468[355] = 42'b100000000000000100100000000000000000001000;
    n1468[354] = 42'b100000000000000010100000000000000000001000;
    n1468[353] = 42'b100000000000001000000000000000000000001010;
    n1468[352] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[351] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[350] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[349] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[348] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[347] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[346] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[345] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[344] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[343] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[342] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[341] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[340] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[339] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[338] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[337] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[336] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[335] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[334] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[333] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[332] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[331] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[330] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[329] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[328] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[327] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[326] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[325] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[324] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[323] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[322] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[321] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[320] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[319] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[318] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[317] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[316] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[315] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[314] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[313] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[312] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[311] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[310] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[309] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[308] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[307] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[306] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[305] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[304] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[303] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[302] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[301] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[300] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[299] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[298] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[297] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[296] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[295] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[294] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[293] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[292] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[291] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[290] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[289] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[288] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[287] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[286] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[285] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[284] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[283] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[282] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[281] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[280] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[279] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[278] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[277] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[276] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[275] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[274] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[273] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[272] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[271] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[270] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[269] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[268] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[267] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[266] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[265] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[264] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[263] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[262] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[261] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[260] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[259] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[258] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[257] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[256] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[255] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[254] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[253] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[252] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[251] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[250] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[249] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[248] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[247] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[246] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[245] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[244] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[243] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[242] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[241] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[240] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[239] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[238] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[237] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[236] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[235] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[234] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[233] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[232] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[231] = 42'b101000011000111000000000000000000000011100;
    n1468[230] = 42'b000001000010010000000000000000000001000000;
    n1468[229] = 42'b000000011000010010000000000000000000000000;
    n1468[228] = 42'b000001000010100000000000000000000001100011;
    n1468[227] = 42'b100000000000000100100000000000000000001000;
    n1468[226] = 42'b100000000000000010100000000000000000001000;
    n1468[225] = 42'b100000000000001000000000000000000000001010;
    n1468[224] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[223] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[222] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[221] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[220] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[219] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[218] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[217] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[216] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[215] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[214] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[213] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[212] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[211] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[210] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[209] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[208] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[207] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[206] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[205] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[204] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[203] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[202] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[201] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[200] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[199] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[198] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[197] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[196] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[195] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[194] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[193] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[192] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[191] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[190] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[189] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[188] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[187] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[186] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[185] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[184] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[183] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[182] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[181] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[180] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[179] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[178] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[177] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[176] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[175] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[174] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[173] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[172] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[171] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[170] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[169] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[168] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[167] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[166] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[165] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[164] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[163] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[162] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[161] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[160] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[159] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[158] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[157] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[156] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[155] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[154] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[153] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[152] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[151] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[150] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[149] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[148] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[147] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[146] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[145] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[144] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[143] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[142] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[141] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[140] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[139] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[138] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[137] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[136] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[135] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[134] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[133] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[132] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[131] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[130] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[129] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[128] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[127] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[126] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[125] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[124] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[123] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[122] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[121] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[120] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[119] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[118] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[117] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[116] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[115] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[114] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[113] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[112] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[111] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[110] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[109] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[108] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[107] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[106] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[105] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[104] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[103] = 42'b101000011100111000000000000000000000011100;
    n1468[102] = 42'b000001000110010000000000000000000001000000;
    n1468[101] = 42'b000000011000010010000000000000000000000000;
    n1468[100] = 42'b000001000010100000000000000000000001100011;
    n1468[99] = 42'b100000000000000100100000000000000000001000;
    n1468[98] = 42'b100000000000000010100000000000000000001000;
    n1468[97] = 42'b100000000000001000000000000000000000001010;
    n1468[96] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[95] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[94] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[93] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[92] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[91] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[90] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[89] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[88] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[87] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[86] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[85] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[84] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[83] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[82] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[81] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[80] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[79] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[78] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[77] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[76] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[75] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[74] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[73] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[72] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[71] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[70] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[69] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[68] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[67] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[66] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[65] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[64] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[63] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[62] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[61] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[60] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[59] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[58] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[57] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[56] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[55] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[54] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[53] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[52] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[51] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[50] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[49] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[48] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[47] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[46] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[45] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[44] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[43] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[42] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[41] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[40] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[39] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[38] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[37] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[36] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[35] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[34] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[33] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[32] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[31] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[30] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[29] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[28] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[27] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[26] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[25] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[24] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[23] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[22] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[21] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[20] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[19] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[18] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[17] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[16] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[15] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[14] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[13] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[12] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[11] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[10] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[9] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[8] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[7] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[6] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[5] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[4] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[3] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[2] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[1] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    n1468[0] = 42'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
    end
  assign n1469_data = n1468[n1423_o];
  /* HUC6280_MC.vhd:6988:54  */
endmodule

module huc6280_cpu
  (input  clk,
   input  rst_n,
   input  ce,
   input  [7:0] di,
   input  rdy,
   input  nmi_n,
   input  irq1_n,
   input  irq2_n,
   input  irqt_n,
   input  vdcnum,
   output [20:0] a_out,
   output [7:0] dout,
   output we_n,
   output mcycle,
   output cs);
  wire en;
  wire [7:0] a;
  wire [7:0] x;
  wire [7:0] y;
  wire [7:0] sp;
  wire [7:0] p;
  wire [15:0] pc;
  wire [15:0] aa;
  wire [7:0] t;
  wire [7:0] dr;
  wire [7:0] sh;
  wire [7:0] dh;
  wire [7:0] lh;
  wire [63:0] mpr;
  wire [7:0] ir;
  wire [4:0] state;
  wire [43:0] mc;
  wire [7:0] next_ir;
  wire [4:0] next_state;
  wire last_cycle;
  wire branch_taken;
  wire mem_inst;
  wire talt;
  wire [15:0] addr_bus;
  wire [7:0] mpr_out;
  wire [7:0] mpr_last;
  wire [6:0] alu_ctrl;
  wire [7:0] alu_l;
  wire [7:0] alu_out;
  wire co;
  wire vo;
  wire no;
  wire zo;
  wire [7:0] mask;
  wire got_int;
  wire res_int;
  wire nmi_int;
  wire irq1_int;
  wire irq2_int;
  wire irqt_int;
  wire brk_int;
  wire old_nmi_n;
  wire nmi_sync;
  wire nmi_active;
  wire n410_o;
  wire n412_o;
  wire [7:0] n413_o;
  wire [7:0] n415_o;
  wire [4:0] n418_o;
  wire n420_o;
  wire n422_o;
  wire n423_o;
  wire [2:0] n424_o;
  wire n425_o;
  wire n426_o;
  wire n428_o;
  wire n429_o;
  wire n431_o;
  wire n432_o;
  wire n433_o;
  wire n435_o;
  wire n436_o;
  wire n438_o;
  wire n439_o;
  wire n440_o;
  wire n442_o;
  wire n443_o;
  wire n445_o;
  wire n446_o;
  wire n447_o;
  wire n449_o;
  wire n450_o;
  wire n452_o;
  wire [7:0] n453_o;
  reg n455_o;
  wire [3:0] n456_o;
  wire n458_o;
  wire n460_o;
  wire n461_o;
  wire [2:0] n462_o;
  wire n466_o;
  wire n467_o;
  wire n470_o;
  wire n472_o;
  wire n473_o;
  wire n478_o;
  wire n480_o;
  wire n481_o;
  wire n483_o;
  wire n484_o;
  wire n486_o;
  wire n487_o;
  wire n489_o;
  wire n490_o;
  wire n492_o;
  wire n493_o;
  wire n495_o;
  wire n496_o;
  wire n498_o;
  wire n499_o;
  wire n501_o;
  wire n502_o;
  wire n504_o;
  wire n505_o;
  wire n507_o;
  wire n508_o;
  wire n510_o;
  wire n511_o;
  wire n513_o;
  wire n514_o;
  wire n516_o;
  wire n517_o;
  wire n519_o;
  wire n520_o;
  wire n522_o;
  wire n523_o;
  wire n525_o;
  wire n526_o;
  wire n528_o;
  wire n529_o;
  wire n531_o;
  wire n532_o;
  wire n534_o;
  wire n535_o;
  wire n537_o;
  wire n538_o;
  wire n540_o;
  wire n541_o;
  wire n543_o;
  wire n544_o;
  wire n546_o;
  wire n547_o;
  wire n549_o;
  wire n550_o;
  wire n552_o;
  wire n553_o;
  wire n555_o;
  wire n556_o;
  wire n558_o;
  wire n559_o;
  wire n561_o;
  wire n562_o;
  wire n564_o;
  wire n565_o;
  wire n567_o;
  wire n568_o;
  wire n570_o;
  wire n571_o;
  wire n573_o;
  wire n574_o;
  wire n576_o;
  wire n577_o;
  wire n579_o;
  wire n580_o;
  wire n582_o;
  wire n583_o;
  wire n584_o;
  wire [1:0] n588_o;
  wire n589_o;
  wire n590_o;
  wire n592_o;
  wire n593_o;
  wire n594_o;
  wire n595_o;
  wire [4:0] n597_o;
  wire [4:0] n599_o;
  wire n601_o;
  wire n602_o;
  wire n603_o;
  wire [4:0] n605_o;
  wire [4:0] n607_o;
  wire n609_o;
  wire [4:0] n611_o;
  wire [4:0] n613_o;
  wire n615_o;
  wire n617_o;
  wire n619_o;
  wire n620_o;
  wire [4:0] n622_o;
  wire [4:0] n624_o;
  wire n626_o;
  wire [3:0] n627_o;
  reg [4:0] n628_o;
  wire n632_o;
  wire n645_o;
  wire n646_o;
  wire n650_o;
  wire n653_o;
  wire n655_o;
  wire n656_o;
  wire n657_o;
  wire n659_o;
  wire [1:0] mcode_m_state_ctrl;
  wire [2:0] mcode_m_addr_bus;
  wire [1:0] mcode_m_load_sdlh;
  wire [2:0] mcode_m_load_p;
  wire [2:0] mcode_m_load_t;
  wire [5:0] mcode_m_addr_ctrl;
  wire [2:0] mcode_m_load_pc;
  wire [2:0] mcode_m_load_sp;
  wire [2:0] mcode_m_axy_ctrl;
  wire [3:0] mcode_m_alubus_ctrl;
  wire [3:0] mcode_m_out_bus;
  wire mcode_m_mem_cycle;
  wire [6:0] mcode_m_alu_ctrl;
  wire [43:0] n665_o;
  wire n671_o;
  wire n673_o;
  wire n675_o;
  wire n676_o;
  wire n677_o;
  wire n679_o;
  wire n681_o;
  wire n683_o;
  wire n684_o;
  wire n685_o;
  wire n686_o;
  wire n687_o;
  wire n688_o;
  wire n689_o;
  wire [4:0] n690_o;
  wire [2:0] n694_o;
  wire n696_o;
  wire n698_o;
  wire n700_o;
  wire n702_o;
  wire n704_o;
  wire n706_o;
  wire n708_o;
  wire [6:0] n709_o;
  reg [7:0] n718_o;
  wire [3:0] n720_o;
  wire n722_o;
  wire n724_o;
  wire n726_o;
  wire n728_o;
  wire n730_o;
  wire n732_o;
  wire n734_o;
  wire n736_o;
  wire n738_o;
  wire n740_o;
  wire n742_o;
  wire [10:0] n744_o;
  reg [7:0] n745_o;
  wire alu_co;
  wire alu_vo;
  wire alu_no;
  wire alu_zo;
  wire [7:0] alu_res;
  wire [2:0] n746_o;
  wire [2:0] n747_o;
  wire n748_o;
  wire n749_o;
  wire n750_o;
  wire n751_o;
  wire n752_o;
  wire n760_o;
  wire n762_o;
  wire n764_o;
  wire n766_o;
  wire n768_o;
  wire n769_o;
  wire n770_o;
  wire n783_o;
  wire [2:0] n785_o;
  wire n787_o;
  wire n789_o;
  wire n791_o;
  wire n793_o;
  wire [3:0] n794_o;
  reg [7:0] n795_o;
  wire n803_o;
  wire [2:0] n805_o;
  wire n807_o;
  wire [7:0] n809_o;
  wire n811_o;
  wire [7:0] n813_o;
  wire n815_o;
  wire [2:0] n816_o;
  reg [7:0] n817_o;
  wire n825_o;
  wire [2:0] n827_o;
  wire n829_o;
  wire n833_o;
  wire n835_o;
  wire [1:0] n836_o;
  wire n837_o;
  wire n839_o;
  wire n840_o;
  wire n842_o;
  wire n845_o;
  wire n846_o;
  wire n848_o;
  wire [3:0] n849_o;
  wire n850_o;
  reg n851_o;
  wire n852_o;
  reg n853_o;
  wire n854_o;
  reg n855_o;
  wire n856_o;
  reg n857_o;
  wire n859_o;
  wire n861_o;
  wire n864_o;
  wire n867_o;
  wire [6:0] n868_o;
  wire n869_o;
  wire n870_o;
  reg n871_o;
  wire n872_o;
  wire n873_o;
  reg n874_o;
  wire n875_o;
  wire n876_o;
  reg n877_o;
  wire n878_o;
  wire n879_o;
  reg n880_o;
  wire n881_o;
  wire n882_o;
  reg n883_o;
  wire n884_o;
  wire n885_o;
  reg n886_o;
  wire n887_o;
  wire n888_o;
  reg n889_o;
  wire n890_o;
  wire n891_o;
  reg n892_o;
  wire n894_o;
  wire n896_o;
  wire n897_o;
  wire n899_o;
  wire [7:0] n900_o;
  wire n908_o;
  wire [1:0] n910_o;
  wire n912_o;
  wire n914_o;
  wire n916_o;
  wire [2:0] n917_o;
  reg [7:0] n918_o;
  reg [7:0] n919_o;
  reg [7:0] n920_o;
  wire n936_o;
  wire n947_o;
  wire n948_o;
  wire n949_o;
  wire [7:0] n950_o;
  wire [7:0] n951_o;
  wire n952_o;
  wire [7:0] n953_o;
  wire [7:0] n954_o;
  wire n955_o;
  wire [7:0] n956_o;
  wire [7:0] n957_o;
  wire n958_o;
  wire [7:0] n959_o;
  wire [7:0] n960_o;
  wire n961_o;
  wire [7:0] n962_o;
  wire [7:0] n963_o;
  wire n964_o;
  wire [7:0] n965_o;
  wire [7:0] n966_o;
  wire n967_o;
  wire [7:0] n968_o;
  wire [7:0] n969_o;
  wire n970_o;
  wire [7:0] n971_o;
  wire [7:0] n972_o;
  wire [63:0] n973_o;
  wire n976_o;
  wire n977_o;
  wire [63:0] n980_o;
  wire [7:0] n984_o;
  wire n985_o;
  wire [7:0] n986_o;
  wire [7:0] n987_o;
  wire n988_o;
  wire [7:0] n989_o;
  wire [7:0] n990_o;
  wire n991_o;
  wire [7:0] n992_o;
  wire [7:0] n993_o;
  wire n994_o;
  wire [7:0] n995_o;
  wire [7:0] n996_o;
  wire n997_o;
  wire [7:0] n998_o;
  wire [7:0] n999_o;
  wire n1000_o;
  wire [7:0] n1001_o;
  wire [7:0] n1002_o;
  wire n1003_o;
  wire [7:0] n1004_o;
  wire [7:0] n1005_o;
  wire n1006_o;
  wire [7:0] n1007_o;
  wire [3:0] n1008_o;
  wire n1010_o;
  wire n1012_o;
  wire n1014_o;
  wire n1016_o;
  wire [2:0] n1017_o;
  wire n1018_o;
  wire [3:0] n1019_o;
  wire [3:0] n1020_o;
  wire [7:0] n1021_o;
  wire n1023_o;
  wire [7:0] n1024_o;
  wire n1026_o;
  wire [7:0] n1027_o;
  wire n1029_o;
  wire [6:0] n1031_o;
  reg [7:0] n1032_o;
  wire [3:0] n1035_o;
  wire n1037_o;
  wire n1038_o;
  wire n1039_o;
  wire n1042_o;
  wire n1047_o;
  wire [15:0] ag_pc;
  wire [15:0] ag_aa;
  wire [2:0] n1054_o;
  wire [5:0] n1055_o;
  wire n1060_o;
  wire n1062_o;
  wire n1063_o;
  wire n1064_o;
  wire n1065_o;
  wire n1066_o;
  wire n1067_o;
  wire n1068_o;
  wire n1070_o;
  wire n1072_o;
  wire n1084_o;
  wire n1086_o;
  wire n1087_o;
  wire n1088_o;
  wire n1089_o;
  wire n1090_o;
  wire n1091_o;
  wire n1092_o;
  wire n1093_o;
  wire n1094_o;
  wire n1095_o;
  wire n1096_o;
  wire n1097_o;
  wire n1099_o;
  wire n1101_o;
  wire n1102_o;
  wire n1103_o;
  wire n1104_o;
  wire n1105_o;
  wire n1106_o;
  wire n1107_o;
  wire n1108_o;
  wire n1109_o;
  wire n1110_o;
  wire n1111_o;
  wire n1112_o;
  wire n1113_o;
  wire n1114_o;
  wire n1122_o;
  wire n1123_o;
  wire n1124_o;
  wire n1125_o;
  wire n1126_o;
  wire n1127_o;
  wire n1128_o;
  wire n1154_o;
  wire n1155_o;
  wire n1156_o;
  wire n1157_o;
  wire [2:0] n1161_o;
  wire n1163_o;
  wire n1165_o;
  wire [15:0] n1167_o;
  wire n1169_o;
  wire [7:0] n1170_o;
  wire [15:0] n1172_o;
  wire n1174_o;
  wire n1176_o;
  wire [3:0] n1178_o;
  wire n1179_o;
  wire [3:0] n1181_o;
  wire n1182_o;
  wire [3:0] n1184_o;
  wire n1185_o;
  wire [3:0] n1187_o;
  wire n1188_o;
  wire [3:0] n1190_o;
  wire n1191_o;
  wire [3:0] n1193_o;
  wire n1194_o;
  wire [3:0] n1196_o;
  wire [3:0] n1197_o;
  wire [3:0] n1198_o;
  wire [3:0] n1199_o;
  wire [3:0] n1200_o;
  wire [3:0] n1201_o;
  wire [3:0] n1202_o;
  wire n1204_o;
  wire [11:0] n1206_o;
  wire [13:0] n1208_o;
  wire [1:0] n1209_o;
  wire n1212_o;
  wire n1215_o;
  wire [1:0] n1217_o;
  reg [1:0] n1218_o;
  wire n1220_o;
  wire [15:0] n1221_o;
  wire n1223_o;
  wire [15:0] n1224_o;
  wire n1226_o;
  wire [7:0] n1227_o;
  wire [1:0] n1228_o;
  wire [1:0] n1229_o;
  wire [1:0] n1230_o;
  wire [1:0] n1231_o;
  wire [1:0] n1232_o;
  wire [1:0] n1233_o;
  wire [1:0] n1234_o;
  wire [1:0] n1235_o;
  reg [1:0] n1236_o;
  wire [1:0] n1237_o;
  wire [1:0] n1238_o;
  wire [1:0] n1239_o;
  wire [1:0] n1240_o;
  wire [1:0] n1241_o;
  wire [1:0] n1242_o;
  wire [1:0] n1243_o;
  wire [1:0] n1244_o;
  wire [1:0] n1245_o;
  reg [1:0] n1246_o;
  wire [11:0] n1247_o;
  wire [11:0] n1248_o;
  wire [11:0] n1249_o;
  wire [11:0] n1250_o;
  wire [11:0] n1251_o;
  wire [11:0] n1252_o;
  wire [11:0] n1253_o;
  wire [11:0] n1254_o;
  reg [11:0] n1255_o;
  wire [12:0] n1257_o;
  wire [2:0] n1259_o;
  wire n1261_o;
  wire [7:0] n1262_o;
  wire [2:0] n1263_o;
  wire [2:0] n1266_o;
  wire n1271_o;
  wire [6:0] n1273_o;
  wire n1275_o;
  wire n1277_o;
  wire n1278_o;
  wire n1279_o;
  wire n1281_o;
  wire n1286_o;
  wire [7:0] n1287_o;
  reg [7:0] n1288_q;
  wire [7:0] n1289_o;
  reg [7:0] n1290_q;
  wire [7:0] n1291_o;
  reg [7:0] n1292_q;
  wire [7:0] n1293_o;
  reg [7:0] n1294_q;
  wire [7:0] n1295_o;
  reg [7:0] n1296_q;
  wire [7:0] n1297_o;
  reg [7:0] n1298_q;
  wire [7:0] n1299_o;
  reg [7:0] n1300_q;
  wire [7:0] n1301_o;
  reg [7:0] n1302_q;
  wire [7:0] n1303_o;
  reg [7:0] n1304_q;
  wire [7:0] n1305_o;
  reg [7:0] n1306_q;
  wire [63:0] n1307_o;
  reg [63:0] n1308_q;
  wire [7:0] n1309_o;
  reg [7:0] n1310_q;
  wire [4:0] n1311_o;
  reg [4:0] n1312_q;
  wire n1313_o;
  reg n1314_q;
  wire [15:0] n1315_o;
  wire n1316_o;
  wire n1317_o;
  wire [7:0] n1318_o;
  reg [7:0] n1319_q;
  wire [6:0] n1320_o;
  wire n1321_o;
  reg n1322_q;
  wire n1323_o;
  reg n1324_q;
  wire n1325_o;
  reg n1326_q;
  wire n1327_o;
  reg n1328_q;
  wire n1329_o;
  reg n1330_q;
  wire n1331_o;
  reg n1332_q;
  wire n1333_o;
  reg n1334_q;
  wire n1335_o;
  reg n1336_q;
  wire n1337_o;
  reg n1338_q;
  wire [20:0] n1339_o;
  wire n1340_o;
  reg n1341_q;
  wire n1342_o;
  wire n1343_o;
  wire n1344_o;
  wire n1345_o;
  wire n1346_o;
  wire n1347_o;
  wire n1348_o;
  wire n1349_o;
  wire [1:0] n1350_o;
  reg n1351_o;
  wire [1:0] n1352_o;
  reg n1353_o;
  wire n1354_o;
  wire n1355_o;
  wire [7:0] n1356_o;
  wire [7:0] n1357_o;
  wire [7:0] n1358_o;
  wire [7:0] n1359_o;
  wire [7:0] n1360_o;
  wire [7:0] n1361_o;
  wire [7:0] n1362_o;
  wire [7:0] n1363_o;
  wire [1:0] n1364_o;
  reg [7:0] n1365_o;
  wire [1:0] n1366_o;
  reg [7:0] n1367_o;
  wire n1368_o;
  wire [7:0] n1369_o;
  assign a_out = n1339_o;
  assign dout = n1032_o;
  assign we_n = n1042_o;
  assign mcycle = n1286_o;
  assign cs = n1341_q;
  /* HUC6280_CPU.vhd:32:16  */
  assign en = n410_o; // (signal)
  /* HUC6280_CPU.vhd:35:16  */
  assign a = n1288_q; // (signal)
  /* HUC6280_CPU.vhd:36:16  */
  assign x = n1290_q; // (signal)
  /* HUC6280_CPU.vhd:37:16  */
  assign y = n1292_q; // (signal)
  /* HUC6280_CPU.vhd:38:16  */
  assign sp = n1294_q; // (signal)
  /* HUC6280_CPU.vhd:39:16  */
  assign p = n1296_q; // (signal)
  /* HUC6280_CPU.vhd:40:16  */
  assign pc = ag_pc; // (signal)
  /* HUC6280_CPU.vhd:41:16  */
  assign aa = ag_aa; // (signal)
  /* HUC6280_CPU.vhd:42:16  */
  assign t = n1298_q; // (signal)
  /* HUC6280_CPU.vhd:43:16  */
  assign dr = n1300_q; // (signal)
  /* HUC6280_CPU.vhd:44:16  */
  assign sh = n1302_q; // (signal)
  /* HUC6280_CPU.vhd:45:16  */
  assign dh = n1304_q; // (signal)
  /* HUC6280_CPU.vhd:46:16  */
  assign lh = n1306_q; // (signal)
  /* HUC6280_CPU.vhd:47:16  */
  assign mpr = n1308_q; // (signal)
  /* HUC6280_CPU.vhd:50:16  */
  assign ir = n1310_q; // (signal)
  /* HUC6280_CPU.vhd:51:16  */
  assign state = n1312_q; // (signal)
  /* HUC6280_CPU.vhd:52:16  */
  assign mc = n665_o; // (signal)
  /* HUC6280_CPU.vhd:53:16  */
  assign next_ir = n413_o; // (signal)
  /* HUC6280_CPU.vhd:54:16  */
  assign next_state = n628_o; // (signal)
  /* HUC6280_CPU.vhd:55:16  */
  assign last_cycle = n646_o; // (signal)
  /* HUC6280_CPU.vhd:56:16  */
  assign branch_taken = n473_o; // (signal)
  /* HUC6280_CPU.vhd:57:16  */
  assign mem_inst = n584_o; // (signal)
  /* HUC6280_CPU.vhd:58:16  */
  assign talt = n1314_q; // (signal)
  /* HUC6280_CPU.vhd:61:16  */
  assign addr_bus = n1315_o; // (signal)
  /* HUC6280_CPU.vhd:62:16  */
  assign mpr_out = n986_o; // (signal)
  /* HUC6280_CPU.vhd:63:16  */
  assign mpr_last = n1319_q; // (signal)
  /* HUC6280_CPU.vhd:66:16  */
  assign alu_ctrl = n1320_o; // (signal)
  /* HUC6280_CPU.vhd:67:16  */
  assign alu_l = n745_o; // (signal)
  /* HUC6280_CPU.vhd:68:16  */
  assign alu_out = alu_res; // (signal)
  /* HUC6280_CPU.vhd:69:16  */
  assign co = alu_co; // (signal)
  /* HUC6280_CPU.vhd:70:16  */
  assign vo = alu_vo; // (signal)
  /* HUC6280_CPU.vhd:71:16  */
  assign no = alu_no; // (signal)
  /* HUC6280_CPU.vhd:72:16  */
  assign zo = alu_zo; // (signal)
  /* HUC6280_CPU.vhd:73:16  */
  assign mask = n718_o; // (signal)
  /* HUC6280_CPU.vhd:76:16  */
  assign got_int = n1322_q; // (signal)
  /* HUC6280_CPU.vhd:77:16  */
  assign res_int = n1324_q; // (signal)
  /* HUC6280_CPU.vhd:78:16  */
  assign nmi_int = n1326_q; // (signal)
  /* HUC6280_CPU.vhd:79:16  */
  assign irq1_int = n1328_q; // (signal)
  /* HUC6280_CPU.vhd:80:16  */
  assign irq2_int = n1330_q; // (signal)
  /* HUC6280_CPU.vhd:81:16  */
  assign irqt_int = n1332_q; // (signal)
  /* HUC6280_CPU.vhd:82:16  */
  assign brk_int = n1157_o; // (signal)
  /* HUC6280_CPU.vhd:83:16  */
  assign old_nmi_n = n1334_q; // (signal)
  /* HUC6280_CPU.vhd:84:16  */
  assign nmi_sync = n1336_q; // (signal)
  /* HUC6280_CPU.vhd:85:16  */
  assign nmi_active = n1338_q; // (signal)
  /* HUC6280_CPU.vhd:89:19  */
  assign n410_o = rdy & ce;
  /* HUC6280_CPU.vhd:91:35  */
  assign n412_o = state != 5'b00000;
  /* HUC6280_CPU.vhd:91:23  */
  assign n413_o = n412_o ? ir : n415_o;
  /* HUC6280_CPU.vhd:91:47  */
  assign n415_o = got_int ? 8'b00000000 : di;
  /* HUC6280_CPU.vhd:99:22  */
  assign n418_o = ir[4:0];
  /* HUC6280_CPU.vhd:99:35  */
  assign n420_o = n418_o == 5'b10000;
  /* HUC6280_CPU.vhd:99:55  */
  assign n422_o = state == 5'b00001;
  /* HUC6280_CPU.vhd:99:45  */
  assign n423_o = n420_o & n422_o;
  /* HUC6280_CPU.vhd:100:32  */
  assign n424_o = ir[7:5];
  /* HUC6280_CPU.vhd:101:68  */
  assign n425_o = p[7];
  /* HUC6280_CPU.vhd:101:63  */
  assign n426_o = ~n425_o;
  /* HUC6280_CPU.vhd:101:33  */
  assign n428_o = n424_o == 3'b000;
  /* HUC6280_CPU.vhd:102:68  */
  assign n429_o = p[7];
  /* HUC6280_CPU.vhd:102:33  */
  assign n431_o = n424_o == 3'b001;
  /* HUC6280_CPU.vhd:103:68  */
  assign n432_o = p[6];
  /* HUC6280_CPU.vhd:103:63  */
  assign n433_o = ~n432_o;
  /* HUC6280_CPU.vhd:103:33  */
  assign n435_o = n424_o == 3'b010;
  /* HUC6280_CPU.vhd:104:68  */
  assign n436_o = p[6];
  /* HUC6280_CPU.vhd:104:33  */
  assign n438_o = n424_o == 3'b011;
  /* HUC6280_CPU.vhd:105:68  */
  assign n439_o = p[0];
  /* HUC6280_CPU.vhd:105:63  */
  assign n440_o = ~n439_o;
  /* HUC6280_CPU.vhd:105:33  */
  assign n442_o = n424_o == 3'b100;
  /* HUC6280_CPU.vhd:106:68  */
  assign n443_o = p[0];
  /* HUC6280_CPU.vhd:106:33  */
  assign n445_o = n424_o == 3'b101;
  /* HUC6280_CPU.vhd:107:68  */
  assign n446_o = p[1];
  /* HUC6280_CPU.vhd:107:63  */
  assign n447_o = ~n446_o;
  /* HUC6280_CPU.vhd:107:33  */
  assign n449_o = n424_o == 3'b110;
  /* HUC6280_CPU.vhd:108:68  */
  assign n450_o = p[1];
  /* HUC6280_CPU.vhd:108:33  */
  assign n452_o = n424_o == 3'b111;
  assign n453_o = {n452_o, n449_o, n445_o, n442_o, n438_o, n435_o, n431_o, n428_o};
  /* HUC6280_CPU.vhd:100:25  */
  always @*
    case (n453_o)
      8'b10000000: n455_o = n450_o;
      8'b01000000: n455_o = n447_o;
      8'b00100000: n455_o = n443_o;
      8'b00010000: n455_o = n440_o;
      8'b00001000: n455_o = n436_o;
      8'b00000100: n455_o = n433_o;
      8'b00000010: n455_o = n429_o;
      8'b00000001: n455_o = n426_o;
      default: n455_o = 1'b0;
    endcase
  /* HUC6280_CPU.vhd:111:25  */
  assign n456_o = ir[3:0];
  /* HUC6280_CPU.vhd:111:38  */
  assign n458_o = n456_o == 4'b1111;
  /* HUC6280_CPU.vhd:111:57  */
  assign n460_o = state == 5'b00101;
  /* HUC6280_CPU.vhd:111:47  */
  assign n461_o = n458_o & n460_o;
  /* HUC6280_CPU.vhd:112:53  */
  assign n462_o = ir[6:4];
  /* HUC6280_CPU.vhd:112:73  */
  assign n466_o = ir[7];
  /* HUC6280_CPU.vhd:112:69  */
  assign n467_o = n1355_o == n466_o;
  /* HUC6280_CPU.vhd:112:25  */
  assign n470_o = n467_o ? 1'b1 : 1'b0;
  /* HUC6280_CPU.vhd:111:17  */
  assign n472_o = n461_o ? n470_o : 1'b0;
  /* HUC6280_CPU.vhd:99:17  */
  assign n473_o = n423_o ? n455_o : n472_o;
  /* HUC6280_CPU.vhd:118:33  */
  assign n478_o = di == 8'b01101001;
  /* HUC6280_CPU.vhd:118:47  */
  assign n480_o = di == 8'b01100101;
  /* HUC6280_CPU.vhd:118:41  */
  assign n481_o = n478_o | n480_o;
  /* HUC6280_CPU.vhd:118:61  */
  assign n483_o = di == 8'b01110101;
  /* HUC6280_CPU.vhd:118:55  */
  assign n484_o = n481_o | n483_o;
  /* HUC6280_CPU.vhd:118:75  */
  assign n486_o = di == 8'b01110010;
  /* HUC6280_CPU.vhd:118:69  */
  assign n487_o = n484_o | n486_o;
  /* HUC6280_CPU.vhd:118:89  */
  assign n489_o = di == 8'b01100001;
  /* HUC6280_CPU.vhd:118:83  */
  assign n490_o = n487_o | n489_o;
  /* HUC6280_CPU.vhd:118:103  */
  assign n492_o = di == 8'b01110001;
  /* HUC6280_CPU.vhd:118:97  */
  assign n493_o = n490_o | n492_o;
  /* HUC6280_CPU.vhd:118:117  */
  assign n495_o = di == 8'b01101101;
  /* HUC6280_CPU.vhd:118:111  */
  assign n496_o = n493_o | n495_o;
  /* HUC6280_CPU.vhd:118:131  */
  assign n498_o = di == 8'b01111101;
  /* HUC6280_CPU.vhd:118:125  */
  assign n499_o = n496_o | n498_o;
  /* HUC6280_CPU.vhd:118:145  */
  assign n501_o = di == 8'b01111001;
  /* HUC6280_CPU.vhd:118:139  */
  assign n502_o = n499_o | n501_o;
  /* HUC6280_CPU.vhd:119:68  */
  assign n504_o = di == 8'b00101001;
  /* HUC6280_CPU.vhd:118:153  */
  assign n505_o = n502_o | n504_o;
  /* HUC6280_CPU.vhd:119:82  */
  assign n507_o = di == 8'b00100101;
  /* HUC6280_CPU.vhd:119:76  */
  assign n508_o = n505_o | n507_o;
  /* HUC6280_CPU.vhd:119:96  */
  assign n510_o = di == 8'b00110101;
  /* HUC6280_CPU.vhd:119:90  */
  assign n511_o = n508_o | n510_o;
  /* HUC6280_CPU.vhd:119:110  */
  assign n513_o = di == 8'b00110010;
  /* HUC6280_CPU.vhd:119:104  */
  assign n514_o = n511_o | n513_o;
  /* HUC6280_CPU.vhd:119:124  */
  assign n516_o = di == 8'b00100001;
  /* HUC6280_CPU.vhd:119:118  */
  assign n517_o = n514_o | n516_o;
  /* HUC6280_CPU.vhd:119:138  */
  assign n519_o = di == 8'b00110001;
  /* HUC6280_CPU.vhd:119:132  */
  assign n520_o = n517_o | n519_o;
  /* HUC6280_CPU.vhd:119:152  */
  assign n522_o = di == 8'b00101101;
  /* HUC6280_CPU.vhd:119:146  */
  assign n523_o = n520_o | n522_o;
  /* HUC6280_CPU.vhd:119:166  */
  assign n525_o = di == 8'b00111101;
  /* HUC6280_CPU.vhd:119:160  */
  assign n526_o = n523_o | n525_o;
  /* HUC6280_CPU.vhd:119:180  */
  assign n528_o = di == 8'b00111001;
  /* HUC6280_CPU.vhd:119:174  */
  assign n529_o = n526_o | n528_o;
  /* HUC6280_CPU.vhd:120:68  */
  assign n531_o = di == 8'b00001001;
  /* HUC6280_CPU.vhd:119:188  */
  assign n532_o = n529_o | n531_o;
  /* HUC6280_CPU.vhd:120:82  */
  assign n534_o = di == 8'b00000101;
  /* HUC6280_CPU.vhd:120:76  */
  assign n535_o = n532_o | n534_o;
  /* HUC6280_CPU.vhd:120:96  */
  assign n537_o = di == 8'b00010101;
  /* HUC6280_CPU.vhd:120:90  */
  assign n538_o = n535_o | n537_o;
  /* HUC6280_CPU.vhd:120:110  */
  assign n540_o = di == 8'b00010010;
  /* HUC6280_CPU.vhd:120:104  */
  assign n541_o = n538_o | n540_o;
  /* HUC6280_CPU.vhd:120:124  */
  assign n543_o = di == 8'b00000001;
  /* HUC6280_CPU.vhd:120:118  */
  assign n544_o = n541_o | n543_o;
  /* HUC6280_CPU.vhd:120:138  */
  assign n546_o = di == 8'b00010001;
  /* HUC6280_CPU.vhd:120:132  */
  assign n547_o = n544_o | n546_o;
  /* HUC6280_CPU.vhd:120:152  */
  assign n549_o = di == 8'b00001101;
  /* HUC6280_CPU.vhd:120:146  */
  assign n550_o = n547_o | n549_o;
  /* HUC6280_CPU.vhd:120:166  */
  assign n552_o = di == 8'b00011101;
  /* HUC6280_CPU.vhd:120:160  */
  assign n553_o = n550_o | n552_o;
  /* HUC6280_CPU.vhd:120:180  */
  assign n555_o = di == 8'b00011001;
  /* HUC6280_CPU.vhd:120:174  */
  assign n556_o = n553_o | n555_o;
  /* HUC6280_CPU.vhd:121:68  */
  assign n558_o = di == 8'b01001001;
  /* HUC6280_CPU.vhd:120:188  */
  assign n559_o = n556_o | n558_o;
  /* HUC6280_CPU.vhd:121:82  */
  assign n561_o = di == 8'b01000101;
  /* HUC6280_CPU.vhd:121:76  */
  assign n562_o = n559_o | n561_o;
  /* HUC6280_CPU.vhd:121:96  */
  assign n564_o = di == 8'b01010101;
  /* HUC6280_CPU.vhd:121:90  */
  assign n565_o = n562_o | n564_o;
  /* HUC6280_CPU.vhd:121:110  */
  assign n567_o = di == 8'b01010010;
  /* HUC6280_CPU.vhd:121:104  */
  assign n568_o = n565_o | n567_o;
  /* HUC6280_CPU.vhd:121:124  */
  assign n570_o = di == 8'b01000001;
  /* HUC6280_CPU.vhd:121:118  */
  assign n571_o = n568_o | n570_o;
  /* HUC6280_CPU.vhd:121:138  */
  assign n573_o = di == 8'b01010001;
  /* HUC6280_CPU.vhd:121:132  */
  assign n574_o = n571_o | n573_o;
  /* HUC6280_CPU.vhd:121:152  */
  assign n576_o = di == 8'b01001101;
  /* HUC6280_CPU.vhd:121:146  */
  assign n577_o = n574_o | n576_o;
  /* HUC6280_CPU.vhd:121:166  */
  assign n579_o = di == 8'b01011101;
  /* HUC6280_CPU.vhd:121:160  */
  assign n580_o = n577_o | n579_o;
  /* HUC6280_CPU.vhd:121:180  */
  assign n582_o = di == 8'b01011001;
  /* HUC6280_CPU.vhd:121:174  */
  assign n583_o = n580_o | n582_o;
  /* HUC6280_CPU.vhd:118:25  */
  assign n584_o = n583_o ? 1'b1 : 1'b0;
  /* HUC6280_CPU.vhd:127:25  */
  assign n588_o = mc[1:0];
  /* HUC6280_CPU.vhd:129:56  */
  assign n589_o = p[5];
  /* HUC6280_CPU.vhd:129:51  */
  assign n590_o = mem_inst & n589_o;
  /* HUC6280_CPU.vhd:129:81  */
  assign n592_o = state == 5'b00000;
  /* HUC6280_CPU.vhd:129:71  */
  assign n593_o = n590_o & n592_o;
  /* HUC6280_CPU.vhd:129:103  */
  assign n594_o = ~got_int;
  /* HUC6280_CPU.vhd:129:91  */
  assign n595_o = n593_o & n594_o;
  /* HUC6280_CPU.vhd:132:61  */
  assign n597_o = state + 5'b00001;
  /* HUC6280_CPU.vhd:129:33  */
  assign n599_o = n595_o ? 5'b01000 : n597_o;
  /* HUC6280_CPU.vhd:128:25  */
  assign n601_o = n588_o == 2'b00;
  /* HUC6280_CPU.vhd:135:37  */
  assign n602_o = p[3];
  /* HUC6280_CPU.vhd:135:46  */
  assign n603_o = ~n602_o;
  /* HUC6280_CPU.vhd:138:61  */
  assign n605_o = state + 5'b00001;
  /* HUC6280_CPU.vhd:135:33  */
  assign n607_o = n603_o ? 5'b00000 : n605_o;
  /* HUC6280_CPU.vhd:134:25  */
  assign n609_o = n588_o == 2'b01;
  /* HUC6280_CPU.vhd:142:61  */
  assign n611_o = state + 5'b00001;
  /* HUC6280_CPU.vhd:141:33  */
  assign n613_o = branch_taken ? n611_o : 5'b00000;
  /* HUC6280_CPU.vhd:140:25  */
  assign n615_o = n588_o == 2'b10;
  /* HUC6280_CPU.vhd:147:38  */
  assign n617_o = a == 8'b00000000;
  /* HUC6280_CPU.vhd:147:53  */
  assign n619_o = lh == 8'b00000000;
  /* HUC6280_CPU.vhd:147:46  */
  assign n620_o = n617_o & n619_o;
  /* HUC6280_CPU.vhd:148:61  */
  assign n622_o = state + 5'b00001;
  /* HUC6280_CPU.vhd:147:33  */
  assign n624_o = n620_o ? n622_o : 5'b01110;
  /* HUC6280_CPU.vhd:146:25  */
  assign n626_o = n588_o == 2'b11;
  assign n627_o = {n626_o, n615_o, n609_o, n601_o};
  /* HUC6280_CPU.vhd:127:17  */
  always @*
    case (n627_o)
      4'b1000: n628_o = n624_o;
      4'b0100: n628_o = n613_o;
      4'b0010: n628_o = n607_o;
      4'b0001: n628_o = n599_o;
      default: n628_o = state;
    endcase
  /* HUC6280_CPU.vhd:160:26  */
  assign n632_o = ~rst_n;
  /* HUC6280_CPU.vhd:171:43  */
  assign n645_o = next_state == 5'b00000;
  /* HUC6280_CPU.vhd:171:27  */
  assign n646_o = n645_o ? 1'b1 : 1'b0;
  /* HUC6280_CPU.vhd:175:26  */
  assign n650_o = ~rst_n;
  /* HUC6280_CPU.vhd:179:42  */
  assign n653_o = state == 5'b01101;
  /* HUC6280_CPU.vhd:181:45  */
  assign n655_o = state == 5'b10011;
  /* HUC6280_CPU.vhd:182:49  */
  assign n656_o = ~talt;
  /* HUC6280_CPU.vhd:181:33  */
  assign n657_o = n655_o ? n656_o : talt;
  /* HUC6280_CPU.vhd:179:33  */
  assign n659_o = n653_o ? 1'b0 : n657_o;
  /* HUC6280_CPU.vhd:188:9  */
  huc6280_mc mcode (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .ir(next_ir),
    .state(next_state),
    .m_state_ctrl(mcode_m_state_ctrl),
    .m_addr_bus(mcode_m_addr_bus),
    .m_load_sdlh(mcode_m_load_sdlh),
    .m_load_p(mcode_m_load_p),
    .m_load_t(mcode_m_load_t),
    .m_addr_ctrl(mcode_m_addr_ctrl),
    .m_load_pc(mcode_m_load_pc),
    .m_load_sp(mcode_m_load_sp),
    .m_axy_ctrl(mcode_m_axy_ctrl),
    .m_alubus_ctrl(mcode_m_alubus_ctrl),
    .m_out_bus(mcode_m_out_bus),
    .m_mem_cycle(mcode_m_mem_cycle),
    .m_alu_ctrl(mcode_m_alu_ctrl));
  assign n665_o = {mcode_m_alu_ctrl, mcode_m_mem_cycle, mcode_m_out_bus, mcode_m_alubus_ctrl, mcode_m_axy_ctrl, mcode_m_load_sp, mcode_m_load_pc, mcode_m_addr_ctrl, mcode_m_load_t, mcode_m_load_p, mcode_m_load_sdlh, mcode_m_addr_bus, mcode_m_state_ctrl};
  /* HUC6280_CPU.vhd:201:23  */
  assign n671_o = ir == 8'b11100011;
  /* HUC6280_CPU.vhd:201:42  */
  assign n673_o = state == 5'b10000;
  /* HUC6280_CPU.vhd:201:56  */
  assign n675_o = state == 5'b10001;
  /* HUC6280_CPU.vhd:201:47  */
  assign n676_o = n673_o | n675_o;
  /* HUC6280_CPU.vhd:201:31  */
  assign n677_o = n671_o & n676_o;
  /* HUC6280_CPU.vhd:203:26  */
  assign n679_o = ir == 8'b11110011;
  /* HUC6280_CPU.vhd:203:45  */
  assign n681_o = state == 5'b01110;
  /* HUC6280_CPU.vhd:203:59  */
  assign n683_o = state == 5'b01111;
  /* HUC6280_CPU.vhd:203:50  */
  assign n684_o = n681_o | n683_o;
  /* HUC6280_CPU.vhd:203:34  */
  assign n685_o = n679_o & n684_o;
  assign n686_o = mc[42];
  /* HUC6280_CPU.vhd:203:17  */
  assign n687_o = n685_o ? talt : n686_o;
  /* HUC6280_CPU.vhd:201:17  */
  assign n688_o = n677_o ? talt : n687_o;
  assign n689_o = mc[43];
  assign n690_o = mc[41:37];
  /* HUC6280_CPU.vhd:210:24  */
  assign n694_o = ir[6:4];
  /* HUC6280_CPU.vhd:211:25  */
  assign n696_o = n694_o == 3'b000;
  /* HUC6280_CPU.vhd:212:25  */
  assign n698_o = n694_o == 3'b001;
  /* HUC6280_CPU.vhd:213:25  */
  assign n700_o = n694_o == 3'b010;
  /* HUC6280_CPU.vhd:214:25  */
  assign n702_o = n694_o == 3'b011;
  /* HUC6280_CPU.vhd:215:25  */
  assign n704_o = n694_o == 3'b100;
  /* HUC6280_CPU.vhd:216:25  */
  assign n706_o = n694_o == 3'b101;
  /* HUC6280_CPU.vhd:217:25  */
  assign n708_o = n694_o == 3'b110;
  assign n709_o = {n708_o, n706_o, n704_o, n702_o, n700_o, n698_o, n696_o};
  /* HUC6280_CPU.vhd:210:17  */
  always @*
    case (n709_o)
      7'b1000000: n718_o = 8'b01000000;
      7'b0100000: n718_o = 8'b00100000;
      7'b0010000: n718_o = 8'b00010000;
      7'b0001000: n718_o = 8'b00001000;
      7'b0000100: n718_o = 8'b00000100;
      7'b0000010: n718_o = 8'b00000010;
      7'b0000001: n718_o = 8'b00000001;
      default: n718_o = 8'b10000000;
    endcase
  /* HUC6280_CPU.vhd:222:17  */
  assign n720_o = mc[31:28];
  /* HUC6280_CPU.vhd:223:41  */
  assign n722_o = n720_o == 4'b0000;
  /* HUC6280_CPU.vhd:224:50  */
  assign n724_o = n720_o == 4'b0001;
  /* HUC6280_CPU.vhd:225:50  */
  assign n726_o = n720_o == 4'b0010;
  /* HUC6280_CPU.vhd:226:50  */
  assign n728_o = n720_o == 4'b0011;
  /* HUC6280_CPU.vhd:227:65  */
  assign n730_o = n720_o == 4'b0100;
  /* HUC6280_CPU.vhd:228:50  */
  assign n732_o = n720_o == 4'b0101;
  /* HUC6280_CPU.vhd:229:50  */
  assign n734_o = n720_o == 4'b1000;
  /* HUC6280_CPU.vhd:230:50  */
  assign n736_o = n720_o == 4'b1001;
  /* HUC6280_CPU.vhd:231:57  */
  assign n738_o = n720_o == 4'b1010;
  /* HUC6280_CPU.vhd:232:57  */
  assign n740_o = n720_o == 4'b1011;
  /* HUC6280_CPU.vhd:233:50  */
  assign n742_o = n720_o == 4'b1100;
  assign n744_o = {n742_o, n740_o, n738_o, n736_o, n734_o, n732_o, n730_o, n728_o, n726_o, n724_o, n722_o};
  /* HUC6280_CPU.vhd:222:9  */
  always @*
    case (n744_o)
      11'b10000000000: n745_o = mask;
      11'b01000000000: n745_o = mpr_out;
      11'b00100000000: n745_o = lh;
      11'b00010000000: n745_o = dh;
      11'b00001000000: n745_o = sh;
      11'b00000100000: n745_o = t;
      11'b00000010000: n745_o = sp;
      11'b00000001000: n745_o = y;
      11'b00000000100: n745_o = x;
      11'b00000000010: n745_o = a;
      11'b00000000001: n745_o = di;
      default: n745_o = 8'b00000000;
    endcase
  /* HUC6280_CPU.vhd:236:9  */
  alu alu (
    .clk(clk),
    .en(en),
    .l(alu_l),
    .r(di),
    .ctrl_fstop(n746_o),
    .ctrl_secop(n747_o),
    .ctrl_fc(n748_o),
    .bcd(n749_o),
    .ci(n750_o),
    .vi(n751_o),
    .ni(n752_o),
    .co(alu_co),
    .vo(alu_vo),
    .no(alu_no),
    .zo(alu_zo),
    .res(alu_res));
  assign n746_o = alu_ctrl[2:0];
  assign n747_o = alu_ctrl[5:3];
  assign n748_o = alu_ctrl[6];
  /* HUC6280_CPU.vhd:243:37  */
  assign n749_o = p[3];
  /* HUC6280_CPU.vhd:244:37  */
  assign n750_o = p[0];
  /* HUC6280_CPU.vhd:245:37  */
  assign n751_o = p[6];
  /* HUC6280_CPU.vhd:246:37  */
  assign n752_o = p[7];
  /* HUC6280_CPU.vhd:257:26  */
  assign n760_o = ~rst_n;
  /* HUC6280_CPU.vhd:263:47  */
  assign n762_o = mc[25];
  /* HUC6280_CPU.vhd:266:47  */
  assign n764_o = mc[26];
  /* HUC6280_CPU.vhd:269:47  */
  assign n766_o = mc[27];
  /* HUC6280_CPU.vhd:262:25  */
  assign n768_o = en & n762_o;
  /* HUC6280_CPU.vhd:262:25  */
  assign n769_o = en & n764_o;
  /* HUC6280_CPU.vhd:262:25  */
  assign n770_o = en & n766_o;
  /* HUC6280_CPU.vhd:278:26  */
  assign n783_o = ~rst_n;
  /* HUC6280_CPU.vhd:282:41  */
  assign n785_o = mc[12:10];
  /* HUC6280_CPU.vhd:283:41  */
  assign n787_o = n785_o == 3'b001;
  /* HUC6280_CPU.vhd:284:41  */
  assign n789_o = n785_o == 3'b010;
  /* HUC6280_CPU.vhd:285:41  */
  assign n791_o = n785_o == 3'b011;
  /* HUC6280_CPU.vhd:286:41  */
  assign n793_o = n785_o == 3'b100;
  assign n794_o = {n793_o, n791_o, n789_o, n787_o};
  /* HUC6280_CPU.vhd:282:33  */
  always @*
    case (n794_o)
      4'b1000: n795_o = di;
      4'b0100: n795_o = y;
      4'b0010: n795_o = x;
      4'b0001: n795_o = alu_out;
      default: n795_o = t;
    endcase
  /* HUC6280_CPU.vhd:295:26  */
  assign n803_o = ~rst_n;
  /* HUC6280_CPU.vhd:299:41  */
  assign n805_o = mc[24:22];
  /* HUC6280_CPU.vhd:300:41  */
  assign n807_o = n805_o == 3'b001;
  /* HUC6280_CPU.vhd:303:85  */
  assign n809_o = sp + 8'b00000001;
  /* HUC6280_CPU.vhd:302:41  */
  assign n811_o = n805_o == 3'b010;
  /* HUC6280_CPU.vhd:305:85  */
  assign n813_o = sp - 8'b00000001;
  /* HUC6280_CPU.vhd:304:41  */
  assign n815_o = n805_o == 3'b011;
  assign n816_o = {n815_o, n811_o, n807_o};
  /* HUC6280_CPU.vhd:299:33  */
  always @*
    case (n816_o)
      3'b100: n817_o = n813_o;
      3'b010: n817_o = n809_o;
      3'b001: n817_o = alu_out;
      default: n817_o = sp;
    endcase
  /* HUC6280_CPU.vhd:315:26  */
  assign n825_o = ~rst_n;
  /* HUC6280_CPU.vhd:319:41  */
  assign n827_o = mc[9:7];
  /* HUC6280_CPU.vhd:320:41  */
  assign n829_o = n827_o == 3'b001;
  /* HUC6280_CPU.vhd:323:41  */
  assign n833_o = n827_o == 3'b010;
  /* HUC6280_CPU.vhd:326:41  */
  assign n835_o = n827_o == 3'b011;
  /* HUC6280_CPU.vhd:329:56  */
  assign n836_o = ir[7:6];
  /* HUC6280_CPU.vhd:330:85  */
  assign n837_o = ir[5];
  /* HUC6280_CPU.vhd:330:57  */
  assign n839_o = n836_o == 2'b00;
  /* HUC6280_CPU.vhd:331:85  */
  assign n840_o = ir[5];
  /* HUC6280_CPU.vhd:331:57  */
  assign n842_o = n836_o == 2'b01;
  /* HUC6280_CPU.vhd:332:57  */
  assign n845_o = n836_o == 2'b10;
  /* HUC6280_CPU.vhd:333:85  */
  assign n846_o = ir[5];
  /* HUC6280_CPU.vhd:333:57  */
  assign n848_o = n836_o == 2'b11;
  assign n849_o = {n848_o, n845_o, n842_o, n839_o};
  assign n850_o = p[0];
  /* HUC6280_CPU.vhd:329:49  */
  always @*
    case (n849_o)
      4'b1000: n851_o = n850_o;
      4'b0100: n851_o = n850_o;
      4'b0010: n851_o = n850_o;
      4'b0001: n851_o = n837_o;
      default: n851_o = n850_o;
    endcase
  assign n852_o = p[2];
  /* HUC6280_CPU.vhd:329:49  */
  always @*
    case (n849_o)
      4'b1000: n853_o = n852_o;
      4'b0100: n853_o = n852_o;
      4'b0010: n853_o = n840_o;
      4'b0001: n853_o = n852_o;
      default: n853_o = n852_o;
    endcase
  assign n854_o = p[3];
  /* HUC6280_CPU.vhd:329:49  */
  always @*
    case (n849_o)
      4'b1000: n855_o = n846_o;
      4'b0100: n855_o = n854_o;
      4'b0010: n855_o = n854_o;
      4'b0001: n855_o = n854_o;
      default: n855_o = n854_o;
    endcase
  assign n856_o = p[6];
  /* HUC6280_CPU.vhd:329:49  */
  always @*
    case (n849_o)
      4'b1000: n857_o = n856_o;
      4'b0100: n857_o = 1'b0;
      4'b0010: n857_o = n856_o;
      4'b0001: n857_o = n856_o;
      default: n857_o = n856_o;
    endcase
  /* HUC6280_CPU.vhd:328:41  */
  assign n859_o = n827_o == 3'b100;
  /* HUC6280_CPU.vhd:336:41  */
  assign n861_o = n827_o == 3'b101;
  /* HUC6280_CPU.vhd:341:41  */
  assign n864_o = n827_o == 3'b110;
  /* HUC6280_CPU.vhd:343:41  */
  assign n867_o = n827_o == 3'b111;
  assign n868_o = {n867_o, n864_o, n861_o, n859_o, n835_o, n833_o, n829_o};
  assign n869_o = di[0];
  assign n870_o = p[0];
  /* HUC6280_CPU.vhd:319:33  */
  always @*
    case (n868_o)
      7'b1000000: n871_o = n870_o;
      7'b0100000: n871_o = n870_o;
      7'b0010000: n871_o = co;
      7'b0001000: n871_o = n851_o;
      7'b0000100: n871_o = n869_o;
      7'b0000010: n871_o = n870_o;
      7'b0000001: n871_o = n870_o;
      default: n871_o = n870_o;
    endcase
  assign n872_o = di[1];
  assign n873_o = p[1];
  /* HUC6280_CPU.vhd:319:33  */
  always @*
    case (n868_o)
      7'b1000000: n874_o = n873_o;
      7'b0100000: n874_o = n873_o;
      7'b0010000: n874_o = zo;
      7'b0001000: n874_o = n873_o;
      7'b0000100: n874_o = n872_o;
      7'b0000010: n874_o = n873_o;
      7'b0000001: n874_o = zo;
      default: n874_o = n873_o;
    endcase
  assign n875_o = di[2];
  assign n876_o = p[2];
  /* HUC6280_CPU.vhd:319:33  */
  always @*
    case (n868_o)
      7'b1000000: n877_o = n876_o;
      7'b0100000: n877_o = n876_o;
      7'b0010000: n877_o = n876_o;
      7'b0001000: n877_o = n853_o;
      7'b0000100: n877_o = n875_o;
      7'b0000010: n877_o = 1'b1;
      7'b0000001: n877_o = n876_o;
      default: n877_o = n876_o;
    endcase
  assign n878_o = di[3];
  assign n879_o = p[3];
  /* HUC6280_CPU.vhd:319:33  */
  always @*
    case (n868_o)
      7'b1000000: n880_o = n879_o;
      7'b0100000: n880_o = n879_o;
      7'b0010000: n880_o = n879_o;
      7'b0001000: n880_o = n855_o;
      7'b0000100: n880_o = n878_o;
      7'b0000010: n880_o = 1'b0;
      7'b0000001: n880_o = n879_o;
      default: n880_o = n879_o;
    endcase
  assign n881_o = di[4];
  assign n882_o = p[4];
  /* HUC6280_CPU.vhd:319:33  */
  always @*
    case (n868_o)
      7'b1000000: n883_o = n882_o;
      7'b0100000: n883_o = n882_o;
      7'b0010000: n883_o = n882_o;
      7'b0001000: n883_o = n882_o;
      7'b0000100: n883_o = n881_o;
      7'b0000010: n883_o = n882_o;
      7'b0000001: n883_o = n882_o;
      default: n883_o = n882_o;
    endcase
  assign n884_o = di[5];
  assign n885_o = p[5];
  /* HUC6280_CPU.vhd:319:33  */
  always @*
    case (n868_o)
      7'b1000000: n886_o = 1'b0;
      7'b0100000: n886_o = 1'b1;
      7'b0010000: n886_o = n885_o;
      7'b0001000: n886_o = n885_o;
      7'b0000100: n886_o = n884_o;
      7'b0000010: n886_o = n885_o;
      7'b0000001: n886_o = n885_o;
      default: n886_o = n885_o;
    endcase
  assign n887_o = di[6];
  assign n888_o = p[6];
  /* HUC6280_CPU.vhd:319:33  */
  always @*
    case (n868_o)
      7'b1000000: n889_o = n888_o;
      7'b0100000: n889_o = n888_o;
      7'b0010000: n889_o = vo;
      7'b0001000: n889_o = n857_o;
      7'b0000100: n889_o = n887_o;
      7'b0000010: n889_o = n888_o;
      7'b0000001: n889_o = n888_o;
      default: n889_o = n888_o;
    endcase
  assign n890_o = di[7];
  assign n891_o = p[7];
  /* HUC6280_CPU.vhd:319:33  */
  always @*
    case (n868_o)
      7'b1000000: n892_o = n891_o;
      7'b0100000: n892_o = n891_o;
      7'b0010000: n892_o = no;
      7'b0001000: n892_o = n891_o;
      7'b0000100: n892_o = n890_o;
      7'b0000010: n892_o = n891_o;
      7'b0000001: n892_o = no;
      default: n892_o = n891_o;
    endcase
  /* HUC6280_CPU.vhd:348:44  */
  assign n894_o = next_ir != 8'b00000000;
  /* HUC6280_CPU.vhd:348:63  */
  assign n896_o = state == 5'b00000;
  /* HUC6280_CPU.vhd:348:53  */
  assign n897_o = n894_o & n896_o;
  /* HUC6280_CPU.vhd:348:33  */
  assign n899_o = n897_o ? 1'b0 : n886_o;
  assign n900_o = {n892_o, n889_o, n899_o, n883_o, n880_o, n877_o, n874_o, n871_o};
  /* HUC6280_CPU.vhd:357:26  */
  assign n908_o = ~rst_n;
  /* HUC6280_CPU.vhd:363:41  */
  assign n910_o = mc[6:5];
  /* HUC6280_CPU.vhd:364:41  */
  assign n912_o = n910_o == 2'b01;
  /* HUC6280_CPU.vhd:365:41  */
  assign n914_o = n910_o == 2'b10;
  /* HUC6280_CPU.vhd:366:41  */
  assign n916_o = n910_o == 2'b11;
  assign n917_o = {n916_o, n914_o, n912_o};
  /* HUC6280_CPU.vhd:363:33  */
  always @*
    case (n917_o)
      3'b100: n918_o = sh;
      3'b010: n918_o = sh;
      3'b001: n918_o = alu_out;
      default: n918_o = sh;
    endcase
  /* HUC6280_CPU.vhd:363:33  */
  always @*
    case (n917_o)
      3'b100: n919_o = dh;
      3'b010: n919_o = alu_out;
      3'b001: n919_o = dh;
      default: n919_o = dh;
    endcase
  /* HUC6280_CPU.vhd:363:33  */
  always @*
    case (n917_o)
      3'b100: n920_o = alu_out;
      3'b010: n920_o = lh;
      3'b001: n920_o = lh;
      default: n920_o = lh;
    endcase
  /* HUC6280_CPU.vhd:375:26  */
  assign n936_o = ~rst_n;
  /* HUC6280_CPU.vhd:386:39  */
  assign n947_o = ir == 8'b01010011;
  /* HUC6280_CPU.vhd:386:47  */
  assign n948_o = n947_o & last_cycle;
  /* HUC6280_CPU.vhd:388:53  */
  assign n949_o = t[0];
  assign n950_o = mpr[63:56];
  /* HUC6280_CPU.vhd:388:49  */
  assign n951_o = n949_o ? a : n950_o;
  /* HUC6280_CPU.vhd:388:53  */
  assign n952_o = t[1];
  assign n953_o = mpr[55:48];
  /* HUC6280_CPU.vhd:388:49  */
  assign n954_o = n952_o ? a : n953_o;
  /* HUC6280_CPU.vhd:388:53  */
  assign n955_o = t[2];
  assign n956_o = mpr[47:40];
  /* HUC6280_CPU.vhd:388:49  */
  assign n957_o = n955_o ? a : n956_o;
  /* HUC6280_CPU.vhd:388:53  */
  assign n958_o = t[3];
  assign n959_o = mpr[39:32];
  /* HUC6280_CPU.vhd:388:49  */
  assign n960_o = n958_o ? a : n959_o;
  /* HUC6280_CPU.vhd:388:53  */
  assign n961_o = t[4];
  assign n962_o = mpr[31:24];
  /* HUC6280_CPU.vhd:388:49  */
  assign n963_o = n961_o ? a : n962_o;
  /* HUC6280_CPU.vhd:388:53  */
  assign n964_o = t[5];
  assign n965_o = mpr[23:16];
  /* HUC6280_CPU.vhd:388:49  */
  assign n966_o = n964_o ? a : n965_o;
  /* HUC6280_CPU.vhd:388:53  */
  assign n967_o = t[6];
  assign n968_o = mpr[15:8];
  /* HUC6280_CPU.vhd:388:49  */
  assign n969_o = n967_o ? a : n968_o;
  /* HUC6280_CPU.vhd:388:53  */
  assign n970_o = t[7];
  assign n971_o = mpr[7:0];
  /* HUC6280_CPU.vhd:388:49  */
  assign n972_o = n970_o ? a : n971_o;
  assign n973_o = {n951_o, n954_o, n957_o, n960_o, n963_o, n966_o, n969_o, n972_o};
  /* HUC6280_CPU.vhd:385:25  */
  assign n976_o = en & n948_o;
  /* HUC6280_CPU.vhd:385:25  */
  assign n977_o = en & n948_o;
  assign n980_o = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
  /* HUC6280_CPU.vhd:398:23  */
  assign n984_o = mpr[63:56];
  /* HUC6280_CPU.vhd:398:33  */
  assign n985_o = t[0];
  /* HUC6280_CPU.vhd:398:27  */
  assign n986_o = n985_o ? n984_o : n989_o;
  /* HUC6280_CPU.vhd:399:38  */
  assign n987_o = mpr[55:48];
  /* HUC6280_CPU.vhd:399:48  */
  assign n988_o = t[1];
  /* HUC6280_CPU.vhd:398:43  */
  assign n989_o = n988_o ? n987_o : n992_o;
  /* HUC6280_CPU.vhd:400:38  */
  assign n990_o = mpr[47:40];
  /* HUC6280_CPU.vhd:400:48  */
  assign n991_o = t[2];
  /* HUC6280_CPU.vhd:399:58  */
  assign n992_o = n991_o ? n990_o : n995_o;
  /* HUC6280_CPU.vhd:401:38  */
  assign n993_o = mpr[39:32];
  /* HUC6280_CPU.vhd:401:48  */
  assign n994_o = t[3];
  /* HUC6280_CPU.vhd:400:58  */
  assign n995_o = n994_o ? n993_o : n998_o;
  /* HUC6280_CPU.vhd:402:38  */
  assign n996_o = mpr[31:24];
  /* HUC6280_CPU.vhd:402:48  */
  assign n997_o = t[4];
  /* HUC6280_CPU.vhd:401:58  */
  assign n998_o = n997_o ? n996_o : n1001_o;
  /* HUC6280_CPU.vhd:403:38  */
  assign n999_o = mpr[23:16];
  /* HUC6280_CPU.vhd:403:48  */
  assign n1000_o = t[5];
  /* HUC6280_CPU.vhd:402:58  */
  assign n1001_o = n1000_o ? n999_o : n1004_o;
  /* HUC6280_CPU.vhd:404:38  */
  assign n1002_o = mpr[15:8];
  /* HUC6280_CPU.vhd:404:48  */
  assign n1003_o = t[6];
  /* HUC6280_CPU.vhd:403:58  */
  assign n1004_o = n1003_o ? n1002_o : n1007_o;
  /* HUC6280_CPU.vhd:405:38  */
  assign n1005_o = mpr[7:0];
  /* HUC6280_CPU.vhd:405:48  */
  assign n1006_o = t[7];
  /* HUC6280_CPU.vhd:404:58  */
  assign n1007_o = n1006_o ? n1005_o : mpr_last;
  /* HUC6280_CPU.vhd:409:17  */
  assign n1008_o = mc[35:32];
  /* HUC6280_CPU.vhd:410:25  */
  assign n1010_o = n1008_o == 4'b0001;
  /* HUC6280_CPU.vhd:411:35  */
  assign n1012_o = n1008_o == 4'b0010;
  /* HUC6280_CPU.vhd:412:35  */
  assign n1014_o = n1008_o == 4'b0011;
  /* HUC6280_CPU.vhd:413:35  */
  assign n1016_o = n1008_o == 4'b0100;
  /* HUC6280_CPU.vhd:414:34  */
  assign n1017_o = p[7:5];
  /* HUC6280_CPU.vhd:414:50  */
  assign n1018_o = ~got_int;
  /* HUC6280_CPU.vhd:414:47  */
  assign n1019_o = {n1017_o, n1018_o};
  /* HUC6280_CPU.vhd:414:66  */
  assign n1020_o = p[3:0];
  /* HUC6280_CPU.vhd:414:63  */
  assign n1021_o = {n1019_o, n1020_o};
  /* HUC6280_CPU.vhd:414:79  */
  assign n1023_o = n1008_o == 4'b0101;
  /* HUC6280_CPU.vhd:415:35  */
  assign n1024_o = pc[15:8];
  /* HUC6280_CPU.vhd:415:49  */
  assign n1026_o = n1008_o == 4'b0110;
  /* HUC6280_CPU.vhd:416:35  */
  assign n1027_o = pc[7:0];
  /* HUC6280_CPU.vhd:416:48  */
  assign n1029_o = n1008_o == 4'b0111;
  assign n1031_o = {n1029_o, n1026_o, n1023_o, n1016_o, n1014_o, n1012_o, n1010_o};
  /* HUC6280_CPU.vhd:409:9  */
  always @*
    case (n1031_o)
      7'b1000000: n1032_o = n1027_o;
      7'b0100000: n1032_o = n1024_o;
      7'b0010000: n1032_o = n1021_o;
      7'b0001000: n1032_o = t;
      7'b0000100: n1032_o = y;
      7'b0000010: n1032_o = x;
      7'b0000001: n1032_o = a;
      default: n1032_o = 8'b00000000;
    endcase
  /* HUC6280_CPU.vhd:422:23  */
  assign n1035_o = mc[35:32];
  /* HUC6280_CPU.vhd:422:31  */
  assign n1037_o = n1035_o != 4'b0000;
  /* HUC6280_CPU.vhd:422:53  */
  assign n1038_o = ~res_int;
  /* HUC6280_CPU.vhd:422:41  */
  assign n1039_o = n1037_o & n1038_o;
  /* HUC6280_CPU.vhd:422:17  */
  assign n1042_o = n1039_o ? 1'b0 : 1'b1;
  /* HUC6280_CPU.vhd:429:26  */
  assign n1047_o = ~rst_n;
  /* HUC6280_CPU.vhd:438:9  */
  huc6280_ag ag (
    .clk(clk),
    .rst_n(rst_n),
    .ce(en),
    .pc_ctrl(n1054_o),
    .addr_ctrl(n1055_o),
    .got_int(got_int),
    .di(di),
    .x(x),
    .y(y),
    .dr(dr),
    .pc(ag_pc),
    .aa(ag_aa));
  /* HUC6280_CPU.vhd:443:39  */
  assign n1054_o = mc[21:19];
  /* HUC6280_CPU.vhd:444:39  */
  assign n1055_o = mc[18:13];
  /* HUC6280_CPU.vhd:457:26  */
  assign n1060_o = ~rst_n;
  /* HUC6280_CPU.vhd:461:36  */
  assign n1062_o = ~res_int;
  /* HUC6280_CPU.vhd:463:42  */
  assign n1063_o = ~nmi_n;
  /* HUC6280_CPU.vhd:463:48  */
  assign n1064_o = n1063_o & old_nmi_n;
  /* HUC6280_CPU.vhd:463:81  */
  assign n1065_o = ~nmi_sync;
  /* HUC6280_CPU.vhd:463:68  */
  assign n1066_o = n1064_o & n1065_o;
  /* HUC6280_CPU.vhd:465:56  */
  assign n1067_o = nmi_active & last_cycle;
  /* HUC6280_CPU.vhd:465:77  */
  assign n1068_o = n1067_o & en;
  /* HUC6280_CPU.vhd:465:33  */
  assign n1070_o = n1068_o ? 1'b0 : nmi_sync;
  /* HUC6280_CPU.vhd:463:33  */
  assign n1072_o = n1066_o ? 1'b1 : n1070_o;
  /* HUC6280_CPU.vhd:474:26  */
  assign n1084_o = ~rst_n;
  /* HUC6280_CPU.vhd:483:38  */
  assign n1086_o = rdy & ce;
  /* HUC6280_CPU.vhd:486:53  */
  assign n1087_o = last_cycle & en;
  /* HUC6280_CPU.vhd:487:52  */
  assign n1088_o = ~got_int;
  /* HUC6280_CPU.vhd:488:62  */
  assign n1089_o = ~irq1_n;
  /* HUC6280_CPU.vhd:488:76  */
  assign n1090_o = ~irq2_n;
  /* HUC6280_CPU.vhd:488:73  */
  assign n1091_o = n1089_o | n1090_o;
  /* HUC6280_CPU.vhd:488:90  */
  assign n1092_o = ~irqt_n;
  /* HUC6280_CPU.vhd:488:87  */
  assign n1093_o = n1091_o | n1092_o;
  /* HUC6280_CPU.vhd:488:111  */
  assign n1094_o = p[2];
  /* HUC6280_CPU.vhd:488:106  */
  assign n1095_o = ~n1094_o;
  /* HUC6280_CPU.vhd:488:102  */
  assign n1096_o = n1093_o & n1095_o;
  /* HUC6280_CPU.vhd:488:121  */
  assign n1097_o = n1096_o | nmi_active;
  /* HUC6280_CPU.vhd:486:33  */
  assign n1099_o = n1122_o ? 1'b0 : nmi_sync;
  /* HUC6280_CPU.vhd:487:41  */
  assign n1101_o = n1088_o ? n1097_o : 1'b0;
  /* HUC6280_CPU.vhd:487:41  */
  assign n1102_o = n1088_o & nmi_active;
  /* HUC6280_CPU.vhd:498:53  */
  assign n1103_o = ~irq1_n;
  /* HUC6280_CPU.vhd:498:73  */
  assign n1104_o = p[2];
  /* HUC6280_CPU.vhd:498:68  */
  assign n1105_o = ~n1104_o;
  /* HUC6280_CPU.vhd:498:64  */
  assign n1106_o = n1103_o & n1105_o;
  /* HUC6280_CPU.vhd:499:53  */
  assign n1107_o = ~irq2_n;
  /* HUC6280_CPU.vhd:499:73  */
  assign n1108_o = p[2];
  /* HUC6280_CPU.vhd:499:68  */
  assign n1109_o = ~n1108_o;
  /* HUC6280_CPU.vhd:499:64  */
  assign n1110_o = n1107_o & n1109_o;
  /* HUC6280_CPU.vhd:500:53  */
  assign n1111_o = ~irqt_n;
  /* HUC6280_CPU.vhd:500:73  */
  assign n1112_o = p[2];
  /* HUC6280_CPU.vhd:500:68  */
  assign n1113_o = ~n1112_o;
  /* HUC6280_CPU.vhd:500:64  */
  assign n1114_o = n1111_o & n1113_o;
  /* HUC6280_CPU.vhd:486:33  */
  assign n1122_o = n1087_o & n1102_o;
  /* HUC6280_CPU.vhd:483:25  */
  assign n1123_o = n1086_o & n1087_o;
  /* HUC6280_CPU.vhd:483:25  */
  assign n1124_o = n1086_o & n1087_o;
  /* HUC6280_CPU.vhd:483:25  */
  assign n1125_o = n1086_o & n1087_o;
  /* HUC6280_CPU.vhd:483:25  */
  assign n1126_o = n1086_o & n1087_o;
  /* HUC6280_CPU.vhd:483:25  */
  assign n1127_o = n1086_o & n1087_o;
  /* HUC6280_CPU.vhd:483:25  */
  assign n1128_o = n1086_o & n1087_o;
  /* HUC6280_CPU.vhd:506:32  */
  assign n1154_o = ir == 8'b00000000;
  /* HUC6280_CPU.vhd:506:52  */
  assign n1155_o = ~got_int;
  /* HUC6280_CPU.vhd:506:40  */
  assign n1156_o = n1154_o & n1155_o;
  /* HUC6280_CPU.vhd:506:24  */
  assign n1157_o = n1156_o ? 1'b1 : 1'b0;
  /* HUC6280_CPU.vhd:511:25  */
  assign n1161_o = mc[4:2];
  /* HUC6280_CPU.vhd:512:25  */
  assign n1163_o = n1161_o == 3'b000;
  /* HUC6280_CPU.vhd:514:25  */
  assign n1165_o = n1161_o == 3'b001;
  /* HUC6280_CPU.vhd:517:51  */
  assign n1167_o = {8'b00100001, sp};
  /* HUC6280_CPU.vhd:516:25  */
  assign n1169_o = n1161_o == 3'b010;
  /* HUC6280_CPU.vhd:519:55  */
  assign n1170_o = aa[7:0];
  /* HUC6280_CPU.vhd:519:51  */
  assign n1172_o = {8'b00100000, n1170_o};
  /* HUC6280_CPU.vhd:518:25  */
  assign n1174_o = n1161_o == 3'b011;
  /* HUC6280_CPU.vhd:523:78  */
  assign n1176_o = state[0];
  /* HUC6280_CPU.vhd:523:71  */
  assign n1178_o = {3'b111, n1176_o};
  /* HUC6280_CPU.vhd:525:78  */
  assign n1179_o = state[0];
  /* HUC6280_CPU.vhd:525:71  */
  assign n1181_o = {3'b110, n1179_o};
  /* HUC6280_CPU.vhd:527:78  */
  assign n1182_o = state[0];
  /* HUC6280_CPU.vhd:527:71  */
  assign n1184_o = {3'b011, n1182_o};
  /* HUC6280_CPU.vhd:529:78  */
  assign n1185_o = state[0];
  /* HUC6280_CPU.vhd:529:71  */
  assign n1187_o = {3'b101, n1185_o};
  /* HUC6280_CPU.vhd:531:78  */
  assign n1188_o = state[0];
  /* HUC6280_CPU.vhd:531:71  */
  assign n1190_o = {3'b100, n1188_o};
  /* HUC6280_CPU.vhd:533:78  */
  assign n1191_o = state[0];
  /* HUC6280_CPU.vhd:533:71  */
  assign n1193_o = {3'b011, n1191_o};
  /* HUC6280_CPU.vhd:535:78  */
  assign n1194_o = state[0];
  /* HUC6280_CPU.vhd:535:71  */
  assign n1196_o = {3'b111, n1194_o};
  /* HUC6280_CPU.vhd:532:33  */
  assign n1197_o = irq2_int ? n1193_o : n1196_o;
  /* HUC6280_CPU.vhd:530:33  */
  assign n1198_o = irq1_int ? n1190_o : n1197_o;
  /* HUC6280_CPU.vhd:528:33  */
  assign n1199_o = irqt_int ? n1187_o : n1198_o;
  /* HUC6280_CPU.vhd:526:33  */
  assign n1200_o = brk_int ? n1184_o : n1199_o;
  /* HUC6280_CPU.vhd:524:33  */
  assign n1201_o = nmi_int ? n1181_o : n1200_o;
  /* HUC6280_CPU.vhd:522:33  */
  assign n1202_o = res_int ? n1178_o : n1201_o;
  /* HUC6280_CPU.vhd:520:25  */
  assign n1204_o = n1161_o == 3'b100;
  /* HUC6280_CPU.vhd:538:72  */
  assign n1206_o = {11'b00000000000, vdcnum};
  /* HUC6280_CPU.vhd:538:81  */
  assign n1208_o = {n1206_o, 2'b00};
  /* HUC6280_CPU.vhd:539:40  */
  assign n1209_o = ir[5:4];
  /* HUC6280_CPU.vhd:540:41  */
  assign n1212_o = n1209_o == 2'b00;
  /* HUC6280_CPU.vhd:541:41  */
  assign n1215_o = n1209_o == 2'b01;
  assign n1217_o = {n1215_o, n1212_o};
  /* HUC6280_CPU.vhd:539:33  */
  always @*
    case (n1217_o)
      2'b10: n1218_o = 2'b10;
      2'b01: n1218_o = 2'b00;
      default: n1218_o = 2'b11;
    endcase
  /* HUC6280_CPU.vhd:537:25  */
  assign n1220_o = n1161_o == 3'b101;
  /* HUC6280_CPU.vhd:545:48  */
  assign n1221_o = {sh, x};
  /* HUC6280_CPU.vhd:544:25  */
  assign n1223_o = n1161_o == 3'b110;
  /* HUC6280_CPU.vhd:547:48  */
  assign n1224_o = {dh, y};
  /* HUC6280_CPU.vhd:546:25  */
  assign n1226_o = n1161_o == 3'b111;
  assign n1227_o = {n1226_o, n1223_o, n1220_o, n1204_o, n1174_o, n1169_o, n1165_o, n1163_o};
  assign n1228_o = pc[1:0];
  assign n1229_o = aa[1:0];
  assign n1230_o = n1167_o[1:0];
  assign n1231_o = n1172_o[1:0];
  assign n1232_o = n1202_o[1:0];
  assign n1233_o = n1221_o[1:0];
  assign n1234_o = n1224_o[1:0];
  assign n1235_o = addr_bus[1:0];
  /* HUC6280_CPU.vhd:511:17  */
  always @*
    case (n1227_o)
      8'b10000000: n1236_o = n1234_o;
      8'b01000000: n1236_o = n1233_o;
      8'b00100000: n1236_o = n1218_o;
      8'b00010000: n1236_o = n1232_o;
      8'b00001000: n1236_o = n1231_o;
      8'b00000100: n1236_o = n1230_o;
      8'b00000010: n1236_o = n1229_o;
      8'b00000001: n1236_o = n1228_o;
      default: n1236_o = n1235_o;
    endcase
  assign n1237_o = pc[3:2];
  assign n1238_o = aa[3:2];
  assign n1239_o = n1167_o[3:2];
  assign n1240_o = n1172_o[3:2];
  assign n1241_o = n1202_o[3:2];
  assign n1242_o = n1208_o[1:0];
  assign n1243_o = n1221_o[3:2];
  assign n1244_o = n1224_o[3:2];
  assign n1245_o = addr_bus[3:2];
  /* HUC6280_CPU.vhd:511:17  */
  always @*
    case (n1227_o)
      8'b10000000: n1246_o = n1244_o;
      8'b01000000: n1246_o = n1243_o;
      8'b00100000: n1246_o = n1242_o;
      8'b00010000: n1246_o = n1241_o;
      8'b00001000: n1246_o = n1240_o;
      8'b00000100: n1246_o = n1239_o;
      8'b00000010: n1246_o = n1238_o;
      8'b00000001: n1246_o = n1237_o;
      default: n1246_o = n1245_o;
    endcase
  assign n1247_o = pc[15:4];
  assign n1248_o = aa[15:4];
  assign n1249_o = n1167_o[15:4];
  assign n1250_o = n1172_o[15:4];
  assign n1251_o = n1208_o[13:2];
  assign n1252_o = n1221_o[15:4];
  assign n1253_o = n1224_o[15:4];
  assign n1254_o = addr_bus[15:4];
  /* HUC6280_CPU.vhd:511:17  */
  always @*
    case (n1227_o)
      8'b10000000: n1255_o = n1253_o;
      8'b01000000: n1255_o = n1252_o;
      8'b00100000: n1255_o = n1251_o;
      8'b00010000: n1255_o = 12'b111111111111;
      8'b00001000: n1255_o = n1250_o;
      8'b00000100: n1255_o = n1249_o;
      8'b00000010: n1255_o = n1248_o;
      8'b00000001: n1255_o = n1247_o;
      default: n1255_o = n1254_o;
    endcase
  /* HUC6280_CPU.vhd:552:39  */
  assign n1257_o = addr_bus[12:0];
  /* HUC6280_CPU.vhd:553:46  */
  assign n1259_o = mc[4:2];
  /* HUC6280_CPU.vhd:553:55  */
  assign n1261_o = n1259_o == 3'b101;
  /* HUC6280_CPU.vhd:553:38  */
  assign n1262_o = n1261_o ? 8'b11111111 : n1369_o;
  /* HUC6280_CPU.vhd:553:100  */
  assign n1263_o = addr_bus[15:13];
  /* HUC6280_CPU.vhd:553:72  */
  assign n1266_o = 3'b111 - n1263_o;
  /* HUC6280_CPU.vhd:557:26  */
  assign n1271_o = ~rst_n;
  /* HUC6280_CPU.vhd:561:38  */
  assign n1273_o = ir[6:0];
  /* HUC6280_CPU.vhd:561:51  */
  assign n1275_o = n1273_o == 7'b1010100;
  /* HUC6280_CPU.vhd:561:73  */
  assign n1277_o = state == 5'b00001;
  /* HUC6280_CPU.vhd:561:63  */
  assign n1278_o = n1275_o & n1277_o;
  /* HUC6280_CPU.vhd:562:49  */
  assign n1279_o = ir[7];
  /* HUC6280_CPU.vhd:560:25  */
  assign n1281_o = en & n1278_o;
  /* HUC6280_CPU.vhd:568:22  */
  assign n1286_o = mc[36];
  /* HUC6280_CPU.vhd:261:17  */
  assign n1287_o = n768_o ? alu_out : a;
  /* HUC6280_CPU.vhd:261:17  */
  always @(posedge clk or posedge n760_o)
    if (n760_o)
      n1288_q <= 8'b00000000;
    else
      n1288_q <= n1287_o;
  /* HUC6280_CPU.vhd:261:17  */
  assign n1289_o = n769_o ? alu_out : x;
  /* HUC6280_CPU.vhd:261:17  */
  always @(posedge clk or posedge n760_o)
    if (n760_o)
      n1290_q <= 8'b00000000;
    else
      n1290_q <= n1289_o;
  /* HUC6280_CPU.vhd:261:17  */
  assign n1291_o = n770_o ? alu_out : y;
  /* HUC6280_CPU.vhd:261:17  */
  always @(posedge clk or posedge n760_o)
    if (n760_o)
      n1292_q <= 8'b00000000;
    else
      n1292_q <= n1291_o;
  /* HUC6280_CPU.vhd:297:17  */
  assign n1293_o = en ? n817_o : sp;
  /* HUC6280_CPU.vhd:297:17  */
  always @(posedge clk or posedge n803_o)
    if (n803_o)
      n1294_q <= 8'b00000000;
    else
      n1294_q <= n1293_o;
  /* HUC6280_CPU.vhd:317:17  */
  assign n1295_o = en ? n900_o : p;
  /* HUC6280_CPU.vhd:317:17  */
  always @(posedge clk or posedge n825_o)
    if (n825_o)
      n1296_q <= 8'b00000100;
    else
      n1296_q <= n1295_o;
  /* HUC6280_CPU.vhd:280:17  */
  assign n1297_o = en ? n795_o : t;
  /* HUC6280_CPU.vhd:280:17  */
  always @(posedge clk or posedge n783_o)
    if (n783_o)
      n1298_q <= 8'b00000000;
    else
      n1298_q <= n1297_o;
  /* HUC6280_CPU.vhd:431:17  */
  assign n1299_o = en ? di : dr;
  /* HUC6280_CPU.vhd:431:17  */
  always @(posedge clk or posedge n1047_o)
    if (n1047_o)
      n1300_q <= 8'b00000000;
    else
      n1300_q <= n1299_o;
  /* HUC6280_CPU.vhd:361:17  */
  assign n1301_o = en ? n918_o : sh;
  /* HUC6280_CPU.vhd:361:17  */
  always @(posedge clk or posedge n908_o)
    if (n908_o)
      n1302_q <= 8'b00000000;
    else
      n1302_q <= n1301_o;
  /* HUC6280_CPU.vhd:361:17  */
  assign n1303_o = en ? n919_o : dh;
  /* HUC6280_CPU.vhd:361:17  */
  always @(posedge clk or posedge n908_o)
    if (n908_o)
      n1304_q <= 8'b00000000;
    else
      n1304_q <= n1303_o;
  /* HUC6280_CPU.vhd:361:17  */
  assign n1305_o = en ? n920_o : lh;
  /* HUC6280_CPU.vhd:361:17  */
  always @(posedge clk or posedge n908_o)
    if (n908_o)
      n1306_q <= 8'b00000000;
    else
      n1306_q <= n1305_o;
  /* HUC6280_CPU.vhd:384:17  */
  assign n1307_o = n976_o ? n973_o : mpr;
  /* HUC6280_CPU.vhd:384:17  */
  always @(posedge clk or posedge n936_o)
    if (n936_o)
      n1308_q <= n980_o;
    else
      n1308_q <= n1307_o;
  /* HUC6280_CPU.vhd:163:17  */
  assign n1309_o = en ? next_ir : ir;
  /* HUC6280_CPU.vhd:163:17  */
  always @(posedge clk or posedge n632_o)
    if (n632_o)
      n1310_q <= 8'b00000000;
    else
      n1310_q <= n1309_o;
  /* HUC6280_CPU.vhd:163:17  */
  assign n1311_o = en ? next_state : state;
  /* HUC6280_CPU.vhd:163:17  */
  always @(posedge clk or posedge n632_o)
    if (n632_o)
      n1312_q <= 5'b00000;
    else
      n1312_q <= n1311_o;
  /* HUC6280_CPU.vhd:177:17  */
  assign n1313_o = en ? n659_o : talt;
  /* HUC6280_CPU.vhd:177:17  */
  always @(posedge clk or posedge n650_o)
    if (n650_o)
      n1314_q <= 1'b0;
    else
      n1314_q <= n1313_o;
  /* HUC6280_CPU.vhd:175:17  */
  assign n1315_o = {n1255_o, n1246_o, n1236_o};
  /* HUC6280_CPU.vhd:373:9  */
  assign n1316_o = ~n936_o;
  /* HUC6280_CPU.vhd:373:9  */
  assign n1317_o = n977_o & n1316_o;
  /* HUC6280_CPU.vhd:384:17  */
  assign n1318_o = n1317_o ? a : mpr_last;
  /* HUC6280_CPU.vhd:384:17  */
  always @(posedge clk)
    n1319_q <= n1318_o;
  /* HUC6280_CPU.vhd:375:17  */
  assign n1320_o = {n689_o, n688_o, n690_o};
  /* HUC6280_CPU.vhd:482:17  */
  assign n1321_o = n1123_o ? n1101_o : got_int;
  /* HUC6280_CPU.vhd:482:17  */
  always @(posedge clk or posedge n1084_o)
    if (n1084_o)
      n1322_q <= 1'b1;
    else
      n1322_q <= n1321_o;
  /* HUC6280_CPU.vhd:482:17  */
  assign n1323_o = n1124_o ? 1'b0 : res_int;
  /* HUC6280_CPU.vhd:482:17  */
  always @(posedge clk or posedge n1084_o)
    if (n1084_o)
      n1324_q <= 1'b1;
    else
      n1324_q <= n1323_o;
  /* HUC6280_CPU.vhd:482:17  */
  assign n1325_o = n1125_o ? nmi_active : nmi_int;
  /* HUC6280_CPU.vhd:482:17  */
  always @(posedge clk or posedge n1084_o)
    if (n1084_o)
      n1326_q <= 1'b0;
    else
      n1326_q <= n1325_o;
  /* HUC6280_CPU.vhd:482:17  */
  assign n1327_o = n1126_o ? n1106_o : irq1_int;
  /* HUC6280_CPU.vhd:482:17  */
  always @(posedge clk or posedge n1084_o)
    if (n1084_o)
      n1328_q <= 1'b0;
    else
      n1328_q <= n1327_o;
  /* HUC6280_CPU.vhd:482:17  */
  assign n1329_o = n1127_o ? n1110_o : irq2_int;
  /* HUC6280_CPU.vhd:482:17  */
  always @(posedge clk or posedge n1084_o)
    if (n1084_o)
      n1330_q <= 1'b0;
    else
      n1330_q <= n1329_o;
  /* HUC6280_CPU.vhd:482:17  */
  assign n1331_o = n1128_o ? n1114_o : irqt_int;
  /* HUC6280_CPU.vhd:482:17  */
  always @(posedge clk or posedge n1084_o)
    if (n1084_o)
      n1332_q <= 1'b0;
    else
      n1332_q <= n1331_o;
  /* HUC6280_CPU.vhd:460:17  */
  assign n1333_o = n1062_o ? nmi_n : old_nmi_n;
  /* HUC6280_CPU.vhd:460:17  */
  always @(posedge clk or posedge n1060_o)
    if (n1060_o)
      n1334_q <= 1'b1;
    else
      n1334_q <= n1333_o;
  /* HUC6280_CPU.vhd:460:17  */
  assign n1335_o = n1062_o ? n1072_o : nmi_sync;
  /* HUC6280_CPU.vhd:460:17  */
  always @(posedge clk or posedge n1060_o)
    if (n1060_o)
      n1336_q <= 1'b0;
    else
      n1336_q <= n1335_o;
  /* HUC6280_CPU.vhd:482:17  */
  assign n1337_o = n1086_o ? n1099_o : nmi_active;
  /* HUC6280_CPU.vhd:482:17  */
  always @(posedge clk or posedge n1084_o)
    if (n1084_o)
      n1338_q <= 1'b0;
    else
      n1338_q <= n1337_o;
  /* HUC6280_CPU.vhd:474:17  */
  assign n1339_o = {n1262_o, n1257_o};
  /* HUC6280_CPU.vhd:559:17  */
  assign n1340_o = n1281_o ? n1279_o : n1341_q;
  /* HUC6280_CPU.vhd:559:17  */
  always @(posedge clk or posedge n1271_o)
    if (n1271_o)
      n1341_q <= 1'b0;
    else
      n1341_q <= n1340_o;
  /* HUC6280_CPU.vhd:451:44  */
  assign n1342_o = dr[0];
  /* HUC6280_CPU.vhd:450:44  */
  assign n1343_o = dr[1];
  /* HUC6280_CPU.vhd:251:36  */
  assign n1344_o = dr[2];
  /* HUC6280_CPU.vhd:250:36  */
  assign n1345_o = dr[3];
  /* HUC6280_CPU.vhd:249:36  */
  assign n1346_o = dr[4];
  /* HUC6280_CPU.vhd:248:28  */
  assign n1347_o = dr[5];
  /* HUC6280_CPU.vhd:247:36  */
  assign n1348_o = dr[6];
  /* HUC6280_CPU.vhd:195:44  */
  assign n1349_o = dr[7];
  /* HUC6280_CPU.vhd:112:30  */
  assign n1350_o = n462_o[1:0];
  /* HUC6280_CPU.vhd:112:30  */
  always @*
    case (n1350_o)
      2'b00: n1351_o = n1342_o;
      2'b01: n1351_o = n1343_o;
      2'b10: n1351_o = n1344_o;
      2'b11: n1351_o = n1345_o;
    endcase
  /* HUC6280_CPU.vhd:112:30  */
  assign n1352_o = n462_o[1:0];
  /* HUC6280_CPU.vhd:112:30  */
  always @*
    case (n1352_o)
      2'b00: n1353_o = n1346_o;
      2'b01: n1353_o = n1347_o;
      2'b10: n1353_o = n1348_o;
      2'b11: n1353_o = n1349_o;
    endcase
  /* HUC6280_CPU.vhd:112:30  */
  assign n1354_o = n462_o[2];
  /* HUC6280_CPU.vhd:112:30  */
  assign n1355_o = n1354_o ? n1353_o : n1351_o;
  /* HUC6280_CPU.vhd:112:30  */
  assign n1356_o = mpr[7:0];
  /* HUC6280_CPU.vhd:112:31  */
  assign n1357_o = mpr[15:8];
  /* HUC6280_CPU.vhd:559:17  */
  assign n1358_o = mpr[23:16];
  /* HUC6280_CPU.vhd:555:9  */
  assign n1359_o = mpr[31:24];
  /* HUC6280_CPU.vhd:553:72  */
  assign n1360_o = mpr[39:32];
  assign n1361_o = mpr[47:40];
  /* HUC6280_CPU.vhd:509:9  */
  assign n1362_o = mpr[55:48];
  assign n1363_o = mpr[63:56];
  /* HUC6280_CPU.vhd:553:71  */
  assign n1364_o = n1266_o[1:0];
  /* HUC6280_CPU.vhd:553:71  */
  always @*
    case (n1364_o)
      2'b00: n1365_o = n1356_o;
      2'b01: n1365_o = n1357_o;
      2'b10: n1365_o = n1358_o;
      2'b11: n1365_o = n1359_o;
    endcase
  /* HUC6280_CPU.vhd:553:71  */
  assign n1366_o = n1266_o[1:0];
  /* HUC6280_CPU.vhd:553:71  */
  always @*
    case (n1366_o)
      2'b00: n1367_o = n1360_o;
      2'b01: n1367_o = n1361_o;
      2'b10: n1367_o = n1362_o;
      2'b11: n1367_o = n1363_o;
    endcase
  /* HUC6280_CPU.vhd:553:71  */
  assign n1368_o = n1266_o[2];
  /* HUC6280_CPU.vhd:553:71  */
  assign n1369_o = n1368_o ? n1367_o : n1365_o;
endmodule

module HUC6280
  (input  CLK,
   input  RST_N,
   input  WAIT_N,
   input  [7:0] DI,
   input  RDY,
   input  NMI_N,
   input  IRQ1_N,
   input  IRQ2_N,
   input  [7:0] K,
   input  VDCNUM,
   output SX,
   output [20:0] A,
   output [7:0] DO,
   output WR_N,
   output RD_N,
   output CE,
   output CEK_N,
   output CE7_N,
   output CER_N,
   output PRE_RD,
   output PRE_WR,
   output HSM,
   output [7:0] O,
   output [23:0] AUD_LDATA,
   output [23:0] AUD_RDATA);
  wire cpu_ce;
  wire cpu_cer;
  wire io_ce;
  wire en;
  wire [7:0] cpu_di;
  wire [7:0] cpu_do;
  wire [20:0] cpu_a;
  wire cpu_we_n;
  wire cpu_cs;
  wire cpu_mcycle;
  wire cpu_irq1_n;
  wire cpu_irq2_n;
  wire cpu_irqt_n;
  wire cpu_rdy;
  wire [4:0] cpu_clk_cnt;
  wire [2:0] io_clk_cnt;
  wire vdc_sel_old;
  wire [7:0] io_buf;
  wire ram_sel;
  wire vdc_sel;
  wire vce_sel;
  wire iop_sel;
  wire psg_sel;
  wire tmr_sel;
  wire int_sel;
  wire io_sel;
  wire [2:0] int_mask;
  wire [9:0] tmr_pre_cnt;
  wire [6:0] tmr_value;
  wire [6:0] tmr_latch;
  wire tmr_en;
  wire tmr_reload;
  wire tmr_irq;
  wire tmr_irq_ack;
  wire n17_o;
  wire n20_o;
  wire n21_o;
  wire n23_o;
  wire n24_o;
  wire n25_o;
  wire n26_o;
  wire n29_o;
  wire n31_o;
  wire n32_o;
  wire n34_o;
  wire n35_o;
  wire n36_o;
  wire n37_o;
  wire n40_o;
  wire [4:0] n42_o;
  wire [4:0] n44_o;
  wire n46_o;
  wire [4:0] n48_o;
  wire n50_o;
  wire n53_o;
  wire [2:0] n56_o;
  wire n58_o;
  wire n61_o;
  wire [2:0] n64_o;
  wire n84_o;
  wire n85_o;
  wire [20:0] core_a_out;
  wire [7:0] core_do;
  wire core_we_n;
  wire core_mcycle;
  wire core_cs;
  wire n91_o;
  wire n92_o;
  wire n93_o;
  wire n94_o;
  wire n95_o;
  wire n96_o;
  wire n97_o;
  wire [5:0] n99_o;
  wire n101_o;
  wire n102_o;
  wire [7:0] n105_o;
  wire n107_o;
  wire [2:0] n108_o;
  wire n110_o;
  wire n111_o;
  wire n112_o;
  wire [7:0] n115_o;
  wire n117_o;
  wire [2:0] n118_o;
  wire n120_o;
  wire n121_o;
  wire n122_o;
  wire n126_o;
  wire n128_o;
  wire n129_o;
  wire n130_o;
  wire n131_o;
  wire n132_o;
  wire n133_o;
  wire n134_o;
  wire n136_o;
  wire n138_o;
  wire n140_o;
  wire n141_o;
  wire n142_o;
  wire n143_o;
  wire n144_o;
  wire n145_o;
  wire n146_o;
  wire n161_o;
  wire n162_o;
  wire n163_o;
  wire n164_o;
  wire n165_o;
  wire n166_o;
  wire n167_o;
  wire n168_o;
  wire [7:0] n170_o;
  wire n172_o;
  wire [2:0] n173_o;
  wire n175_o;
  wire n176_o;
  wire n177_o;
  wire n181_o;
  wire n183_o;
  wire n184_o;
  wire n186_o;
  wire [7:0] n192_o;
  wire n194_o;
  wire [2:0] n195_o;
  wire n197_o;
  wire n198_o;
  wire n199_o;
  wire n203_o;
  wire n205_o;
  wire n206_o;
  wire [1:0] n207_o;
  wire [2:0] n208_o;
  wire n210_o;
  wire n212_o;
  wire [1:0] n213_o;
  reg [2:0] n214_o;
  reg n217_o;
  wire [1:0] n218_o;
  wire n220_o;
  reg n223_o;
  wire n225_o;
  wire n226_o;
  wire n228_o;
  wire [7:0] n238_o;
  wire n240_o;
  wire [2:0] n241_o;
  wire n243_o;
  wire n244_o;
  wire n245_o;
  wire n249_o;
  wire n251_o;
  wire n252_o;
  wire n253_o;
  wire n254_o;
  wire n255_o;
  wire [6:0] n256_o;
  wire n257_o;
  wire n258_o;
  wire n259_o;
  wire n260_o;
  wire [9:0] n262_o;
  wire [6:0] n263_o;
  wire [9:0] n264_o;
  wire [6:0] n265_o;
  wire n267_o;
  wire [9:0] n268_o;
  wire [6:0] n269_o;
  wire n270_o;
  wire n273_o;
  wire [9:0] n275_o;
  wire n277_o;
  wire [6:0] n279_o;
  wire n281_o;
  wire n284_o;
  wire n286_o;
  wire [6:0] n287_o;
  wire n289_o;
  wire n290_o;
  wire [9:0] n291_o;
  wire n292_o;
  wire n294_o;
  wire n296_o;
  wire [6:0] n297_o;
  wire n298_o;
  wire [6:0] n299_o;
  wire n301_o;
  wire [7:0] n322_o;
  wire n324_o;
  wire [2:0] n325_o;
  wire n327_o;
  wire n328_o;
  wire n329_o;
  wire n331_o;
  wire n332_o;
  wire n333_o;
  wire n336_o;
  wire n338_o;
  wire [7:0] n339_o;
  wire n341_o;
  wire n349_o;
  wire [1:0] n350_o;
  wire [4:0] n351_o;
  wire [7:0] n352_o;
  wire n354_o;
  wire [4:0] n355_o;
  wire [5:0] n356_o;
  wire n357_o;
  wire [6:0] n358_o;
  wire n359_o;
  wire [7:0] n360_o;
  wire n362_o;
  wire [1:0] n363_o;
  reg [7:0] n364_o;
  wire n365_o;
  wire [7:0] n366_o;
  wire [7:0] n367_o;
  wire [7:0] n368_o;
  wire [7:0] n369_o;
  wire [7:0] n371_o;
  wire [7:0] n372_o;
  reg n375_q;
  reg n376_q;
  reg n377_q;
  reg [7:0] n378_q;
  reg n379_q;
  reg [4:0] n380_q;
  reg [2:0] n381_q;
  wire n382_o;
  reg n383_q;
  wire [7:0] n384_o;
  reg [7:0] n385_q;
  wire [2:0] n386_o;
  reg [2:0] n387_q;
  reg [9:0] n388_q;
  reg [6:0] n389_q;
  wire [6:0] n390_o;
  reg [6:0] n391_q;
  wire n392_o;
  reg n393_q;
  wire n394_o;
  reg n395_q;
  reg n396_q;
  reg n397_q;
  reg n398_q;
  reg n399_q;
  reg n400_q;
  wire [7:0] n401_o;
  reg [7:0] n402_q;
  localparam [23:0] n403_o = 24'bZ;
  localparam [23:0] n404_o = 24'bZ;
  assign SX = n398_q;
  assign A = cpu_a;
  assign DO = cpu_do;
  assign WR_N = n399_q;
  assign RD_N = n400_q;
  assign CE = n84_o;
  assign CEK_N = n168_o;
  assign CE7_N = n167_o;
  assign CER_N = n166_o;
  assign PRE_RD = n162_o;
  assign PRE_WR = n165_o;
  assign HSM = cpu_cs;
  assign O = n402_q;
  assign AUD_LDATA = n403_o;
  assign AUD_RDATA = n404_o;
  /* HUC6280.vhd:45:16  */
  assign cpu_ce = n375_q; // (signal)
  /* HUC6280.vhd:46:16  */
  assign cpu_cer = n376_q; // (signal)
  /* HUC6280.vhd:47:16  */
  assign io_ce = n377_q; // (signal)
  /* HUC6280.vhd:48:16  */
  assign en = n85_o; // (signal)
  /* HUC6280.vhd:50:16  */
  assign cpu_di = n378_q; // (signal)
  /* HUC6280.vhd:51:16  */
  assign cpu_do = core_do; // (signal)
  /* HUC6280.vhd:52:16  */
  assign cpu_a = core_a_out; // (signal)
  /* HUC6280.vhd:53:16  */
  assign cpu_we_n = core_we_n; // (signal)
  /* HUC6280.vhd:54:16  */
  assign cpu_cs = core_cs; // (signal)
  /* HUC6280.vhd:55:16  */
  assign cpu_mcycle = core_mcycle; // (signal)
  /* HUC6280.vhd:56:16  */
  assign cpu_irq1_n = n92_o; // (signal)
  /* HUC6280.vhd:57:16  */
  assign cpu_irq2_n = n94_o; // (signal)
  /* HUC6280.vhd:58:16  */
  assign cpu_irqt_n = n97_o; // (signal)
  /* HUC6280.vhd:59:16  */
  assign cpu_rdy = n379_q; // (signal)
  /* HUC6280.vhd:61:16  */
  assign cpu_clk_cnt = n380_q; // (signal)
  /* HUC6280.vhd:62:16  */
  assign io_clk_cnt = n381_q; // (signal)
  /* HUC6280.vhd:63:16  */
  assign vdc_sel_old = n383_q; // (signal)
  /* HUC6280.vhd:66:16  */
  assign io_buf = n385_q; // (signal)
  /* HUC6280.vhd:67:16  */
  assign ram_sel = n102_o; // (signal)
  /* HUC6280.vhd:68:16  */
  assign vdc_sel = n112_o; // (signal)
  /* HUC6280.vhd:69:16  */
  assign vce_sel = n122_o; // (signal)
  /* HUC6280.vhd:70:16  */
  assign iop_sel = n177_o; // (signal)
  /* HUC6280.vhd:71:16  */
  assign psg_sel = n329_o; // (signal)
  /* HUC6280.vhd:72:16  */
  assign tmr_sel = n245_o; // (signal)
  /* HUC6280.vhd:73:16  */
  assign int_sel = n199_o; // (signal)
  /* HUC6280.vhd:74:16  */
  assign io_sel = n333_o; // (signal)
  /* HUC6280.vhd:76:16  */
  assign int_mask = n387_q; // (signal)
  /* HUC6280.vhd:77:16  */
  assign tmr_pre_cnt = n388_q; // (signal)
  /* HUC6280.vhd:78:16  */
  assign tmr_value = n389_q; // (signal)
  /* HUC6280.vhd:79:16  */
  assign tmr_latch = n391_q; // (signal)
  /* HUC6280.vhd:80:16  */
  assign tmr_en = n393_q; // (signal)
  /* HUC6280.vhd:81:16  */
  assign tmr_reload = n395_q; // (signal)
  /* HUC6280.vhd:82:16  */
  assign tmr_irq = n396_q; // (signal)
  /* HUC6280.vhd:83:16  */
  assign tmr_irq_ack = n397_q; // (signal)
  /* HUC6280.vhd:90:26  */
  assign n17_o = ~RST_N;
  /* HUC6280.vhd:99:41  */
  assign n20_o = cpu_clk_cnt == 5'b00010;
  /* HUC6280.vhd:99:45  */
  assign n21_o = n20_o & cpu_cs;
  /* HUC6280.vhd:99:79  */
  assign n23_o = cpu_clk_cnt == 5'b01011;
  /* HUC6280.vhd:99:95  */
  assign n24_o = ~cpu_cs;
  /* HUC6280.vhd:99:84  */
  assign n25_o = n23_o & n24_o;
  /* HUC6280.vhd:99:63  */
  assign n26_o = n21_o | n25_o;
  /* HUC6280.vhd:99:25  */
  assign n29_o = n26_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:104:41  */
  assign n31_o = cpu_clk_cnt == 5'b00101;
  /* HUC6280.vhd:104:45  */
  assign n32_o = n31_o & cpu_cs;
  /* HUC6280.vhd:104:79  */
  assign n34_o = cpu_clk_cnt == 5'b10111;
  /* HUC6280.vhd:104:95  */
  assign n35_o = ~cpu_cs;
  /* HUC6280.vhd:104:84  */
  assign n36_o = n34_o & n35_o;
  /* HUC6280.vhd:104:63  */
  assign n37_o = n32_o | n36_o;
  /* HUC6280.vhd:105:33  */
  assign n40_o = WAIT_N ? 1'b1 : 1'b0;
  /* HUC6280.vhd:105:33  */
  assign n42_o = WAIT_N ? 5'b00000 : cpu_clk_cnt;
  /* HUC6280.vhd:110:60  */
  assign n44_o = cpu_clk_cnt + 5'b00001;
  /* HUC6280.vhd:104:25  */
  assign n46_o = n37_o ? n40_o : 1'b0;
  /* HUC6280.vhd:104:25  */
  assign n48_o = n37_o ? n42_o : n44_o;
  /* HUC6280.vhd:114:40  */
  assign n50_o = cpu_clk_cnt == 5'b00001;
  /* HUC6280.vhd:114:25  */
  assign n53_o = n50_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:119:50  */
  assign n56_o = io_clk_cnt + 3'b001;
  /* HUC6280.vhd:120:39  */
  assign n58_o = io_clk_cnt == 3'b101;
  /* HUC6280.vhd:120:25  */
  assign n61_o = n58_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:120:25  */
  assign n64_o = n58_o ? 3'b000 : n56_o;
  /* HUC6280.vhd:127:22  */
  assign n84_o = cpu_ce & cpu_rdy;
  /* HUC6280.vhd:129:22  */
  assign n85_o = cpu_ce & cpu_rdy;
  /* HUC6280.vhd:132:9  */
  huc6280_cpu core (
    .clk(CLK),
    .rst_n(RST_N),
    .ce(cpu_ce),
    .di(cpu_di),
    .rdy(cpu_rdy),
    .nmi_n(NMI_N),
    .irq1_n(cpu_irq1_n),
    .irq2_n(cpu_irq2_n),
    .irqt_n(cpu_irqt_n),
    .vdcnum(VDCNUM),
    .a_out(core_a_out),
    .dout(core_do),
    .we_n(core_we_n),
    .mcycle(core_mcycle),
    .cs(core_cs));
  /* HUC6280.vhd:152:41  */
  assign n91_o = int_mask[1];
  /* HUC6280.vhd:152:30  */
  assign n92_o = IRQ1_N | n91_o;
  /* HUC6280.vhd:153:41  */
  assign n93_o = int_mask[0];
  /* HUC6280.vhd:153:30  */
  assign n94_o = IRQ2_N | n93_o;
  /* HUC6280.vhd:154:23  */
  assign n95_o = ~tmr_irq;
  /* HUC6280.vhd:154:46  */
  assign n96_o = int_mask[2];
  /* HUC6280.vhd:154:35  */
  assign n97_o = n95_o | n96_o;
  /* HUC6280.vhd:156:34  */
  assign n99_o = cpu_a[20:15];
  /* HUC6280.vhd:156:49  */
  assign n101_o = n99_o == 6'b111110;
  /* HUC6280.vhd:156:24  */
  assign n102_o = n101_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:157:34  */
  assign n105_o = cpu_a[20:13];
  /* HUC6280.vhd:157:49  */
  assign n107_o = n105_o == 8'b11111111;
  /* HUC6280.vhd:157:66  */
  assign n108_o = cpu_a[12:10];
  /* HUC6280.vhd:157:81  */
  assign n110_o = n108_o == 3'b000;
  /* HUC6280.vhd:157:57  */
  assign n111_o = n107_o & n110_o;
  /* HUC6280.vhd:157:24  */
  assign n112_o = n111_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:158:34  */
  assign n115_o = cpu_a[20:13];
  /* HUC6280.vhd:158:49  */
  assign n117_o = n115_o == 8'b11111111;
  /* HUC6280.vhd:158:66  */
  assign n118_o = cpu_a[12:10];
  /* HUC6280.vhd:158:81  */
  assign n120_o = n118_o == 3'b001;
  /* HUC6280.vhd:158:57  */
  assign n121_o = n117_o & n120_o;
  /* HUC6280.vhd:158:24  */
  assign n122_o = n121_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:162:26  */
  assign n126_o = ~RST_N;
  /* HUC6280.vhd:171:49  */
  assign n128_o = ~cpu_we_n;
  /* HUC6280.vhd:169:33  */
  assign n129_o = cpu_mcycle ? cpu_we_n : n399_q;
  /* HUC6280.vhd:169:33  */
  assign n130_o = cpu_mcycle ? n128_o : n400_q;
  /* HUC6280.vhd:174:56  */
  assign n131_o = vdc_sel | vce_sel;
  /* HUC6280.vhd:175:51  */
  assign n132_o = vdc_sel | vce_sel;
  /* HUC6280.vhd:175:85  */
  assign n133_o = ~vdc_sel_old;
  /* HUC6280.vhd:175:69  */
  assign n134_o = n132_o & n133_o;
  /* HUC6280.vhd:175:33  */
  assign n136_o = n134_o ? 1'b0 : cpu_rdy;
  /* HUC6280.vhd:178:25  */
  assign n138_o = n141_o ? 1'b1 : n399_q;
  /* HUC6280.vhd:178:25  */
  assign n140_o = n142_o ? 1'b1 : n400_q;
  /* HUC6280.vhd:178:25  */
  assign n141_o = cpu_ce & cpu_rdy;
  /* HUC6280.vhd:178:25  */
  assign n142_o = cpu_ce & cpu_rdy;
  /* HUC6280.vhd:178:25  */
  assign n143_o = cpu_ce ? RDY : cpu_rdy;
  /* HUC6280.vhd:168:25  */
  assign n144_o = cpu_cer ? n129_o : n138_o;
  /* HUC6280.vhd:168:25  */
  assign n145_o = cpu_cer ? n130_o : n140_o;
  /* HUC6280.vhd:168:25  */
  assign n146_o = cpu_cer ? n136_o : n143_o;
  /* HUC6280.vhd:188:28  */
  assign n161_o = cpu_we_n & cpu_mcycle;
  /* HUC6280.vhd:188:43  */
  assign n162_o = n161_o & RST_N;
  /* HUC6280.vhd:189:19  */
  assign n163_o = ~cpu_we_n;
  /* HUC6280.vhd:189:32  */
  assign n164_o = n163_o & cpu_mcycle;
  /* HUC6280.vhd:189:47  */
  assign n165_o = n164_o & RST_N;
  /* HUC6280.vhd:193:18  */
  assign n166_o = ~ram_sel;
  /* HUC6280.vhd:194:18  */
  assign n167_o = ~vdc_sel;
  /* HUC6280.vhd:195:18  */
  assign n168_o = ~vce_sel;
  /* HUC6280.vhd:201:34  */
  assign n170_o = cpu_a[20:13];
  /* HUC6280.vhd:201:49  */
  assign n172_o = n170_o == 8'b11111111;
  /* HUC6280.vhd:201:66  */
  assign n173_o = cpu_a[12:10];
  /* HUC6280.vhd:201:81  */
  assign n175_o = n173_o == 3'b100;
  /* HUC6280.vhd:201:57  */
  assign n176_o = n172_o & n175_o;
  /* HUC6280.vhd:201:24  */
  assign n177_o = n176_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:204:26  */
  assign n181_o = ~RST_N;
  /* HUC6280.vhd:208:63  */
  assign n183_o = ~cpu_we_n;
  /* HUC6280.vhd:208:50  */
  assign n184_o = iop_sel & n183_o;
  /* HUC6280.vhd:207:25  */
  assign n186_o = en & n184_o;
  /* HUC6280.vhd:216:34  */
  assign n192_o = cpu_a[20:13];
  /* HUC6280.vhd:216:49  */
  assign n194_o = n192_o == 8'b11111111;
  /* HUC6280.vhd:216:66  */
  assign n195_o = cpu_a[12:10];
  /* HUC6280.vhd:216:81  */
  assign n197_o = n195_o == 3'b101;
  /* HUC6280.vhd:216:57  */
  assign n198_o = n194_o & n197_o;
  /* HUC6280.vhd:216:24  */
  assign n199_o = n198_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:219:26  */
  assign n203_o = ~RST_N;
  /* HUC6280.vhd:224:42  */
  assign n205_o = int_sel & cpu_cer;
  /* HUC6280.vhd:225:45  */
  assign n206_o = ~cpu_we_n;
  /* HUC6280.vhd:226:51  */
  assign n207_o = cpu_a[1:0];
  /* HUC6280.vhd:228:75  */
  assign n208_o = cpu_do[2:0];
  /* HUC6280.vhd:227:49  */
  assign n210_o = n207_o == 2'b10;
  /* HUC6280.vhd:229:49  */
  assign n212_o = n207_o == 2'b11;
  assign n213_o = {n212_o, n210_o};
  /* HUC6280.vhd:226:41  */
  always @*
    case (n213_o)
      2'b10: n214_o = int_mask;
      2'b01: n214_o = n208_o;
      default: n214_o = int_mask;
    endcase
  /* HUC6280.vhd:226:41  */
  always @*
    case (n213_o)
      2'b10: n217_o = 1'b1;
      2'b01: n217_o = 1'b0;
      default: n217_o = 1'b0;
    endcase
  /* HUC6280.vhd:234:51  */
  assign n218_o = cpu_a[1:0];
  /* HUC6280.vhd:235:49  */
  assign n220_o = n218_o == 2'b10;
  /* HUC6280.vhd:234:41  */
  always @*
    case (n220_o)
      1'b1: n223_o = 1'b1;
      default: n223_o = 1'b0;
    endcase
  /* HUC6280.vhd:225:33  */
  assign n225_o = n206_o ? n217_o : n223_o;
  /* HUC6280.vhd:224:25  */
  assign n226_o = n205_o & n206_o;
  /* HUC6280.vhd:224:25  */
  assign n228_o = n205_o ? n225_o : 1'b0;
  /* HUC6280.vhd:246:34  */
  assign n238_o = cpu_a[20:13];
  /* HUC6280.vhd:246:49  */
  assign n240_o = n238_o == 8'b11111111;
  /* HUC6280.vhd:246:66  */
  assign n241_o = cpu_a[12:10];
  /* HUC6280.vhd:246:81  */
  assign n243_o = n241_o == 3'b011;
  /* HUC6280.vhd:246:57  */
  assign n244_o = n240_o & n243_o;
  /* HUC6280.vhd:246:24  */
  assign n245_o = n244_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:249:26  */
  assign n249_o = ~RST_N;
  /* HUC6280.vhd:257:55  */
  assign n251_o = ~cpu_we_n;
  /* HUC6280.vhd:257:42  */
  assign n252_o = tmr_sel & n251_o;
  /* HUC6280.vhd:257:61  */
  assign n253_o = n252_o & cpu_cer;
  /* HUC6280.vhd:258:41  */
  assign n254_o = cpu_a[0];
  /* HUC6280.vhd:258:45  */
  assign n255_o = ~n254_o;
  /* HUC6280.vhd:260:60  */
  assign n256_o = cpu_do[6:0];
  /* HUC6280.vhd:263:57  */
  assign n257_o = cpu_do[0];
  /* HUC6280.vhd:264:51  */
  assign n258_o = ~tmr_en;
  /* HUC6280.vhd:264:67  */
  assign n259_o = cpu_do[0];
  /* HUC6280.vhd:264:57  */
  assign n260_o = n258_o & n259_o;
  /* HUC6280.vhd:264:41  */
  assign n262_o = n260_o ? 10'b1111111111 : tmr_pre_cnt;
  /* HUC6280.vhd:264:41  */
  assign n263_o = n260_o ? tmr_latch : tmr_value;
  /* HUC6280.vhd:258:33  */
  assign n264_o = n255_o ? tmr_pre_cnt : n262_o;
  /* HUC6280.vhd:258:33  */
  assign n265_o = n255_o ? tmr_value : n263_o;
  /* HUC6280.vhd:258:33  */
  assign n267_o = n255_o ? tmr_en : n257_o;
  /* HUC6280.vhd:257:25  */
  assign n268_o = n253_o ? n264_o : tmr_pre_cnt;
  /* HUC6280.vhd:257:25  */
  assign n269_o = n253_o ? n265_o : tmr_value;
  /* HUC6280.vhd:257:25  */
  assign n270_o = n253_o & n255_o;
  /* HUC6280.vhd:271:25  */
  assign n273_o = tmr_irq_ack ? 1'b0 : tmr_irq;
  /* HUC6280.vhd:278:68  */
  assign n275_o = tmr_pre_cnt - 10'b0000000001;
  /* HUC6280.vhd:279:56  */
  assign n277_o = tmr_pre_cnt == 10'b0000000000;
  /* HUC6280.vhd:280:100  */
  assign n279_o = tmr_value - 7'b0000001;
  /* HUC6280.vhd:281:62  */
  assign n281_o = tmr_value == 7'b0000000;
  /* HUC6280.vhd:281:49  */
  assign n284_o = n281_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:275:25  */
  assign n286_o = n301_o ? 1'b1 : n273_o;
  /* HUC6280.vhd:277:33  */
  assign n287_o = n292_o ? n279_o : n269_o;
  /* HUC6280.vhd:279:41  */
  assign n289_o = n277_o ? n284_o : 1'b0;
  /* HUC6280.vhd:279:41  */
  assign n290_o = n277_o & n281_o;
  /* HUC6280.vhd:275:25  */
  assign n291_o = n298_o ? n275_o : n268_o;
  /* HUC6280.vhd:277:33  */
  assign n292_o = tmr_en & n277_o;
  /* HUC6280.vhd:277:33  */
  assign n294_o = tmr_en ? n289_o : 1'b0;
  /* HUC6280.vhd:277:33  */
  assign n296_o = tmr_en & n290_o;
  /* HUC6280.vhd:288:33  */
  assign n297_o = tmr_reload ? tmr_latch : n287_o;
  /* HUC6280.vhd:275:25  */
  assign n298_o = io_ce & tmr_en;
  /* HUC6280.vhd:275:25  */
  assign n299_o = io_ce ? n297_o : n269_o;
  /* HUC6280.vhd:275:25  */
  assign n301_o = io_ce & n296_o;
  /* HUC6280.vhd:296:34  */
  assign n322_o = cpu_a[20:13];
  /* HUC6280.vhd:296:49  */
  assign n324_o = n322_o == 8'b11111111;
  /* HUC6280.vhd:296:66  */
  assign n325_o = cpu_a[12:10];
  /* HUC6280.vhd:296:81  */
  assign n327_o = n325_o == 3'b010;
  /* HUC6280.vhd:296:57  */
  assign n328_o = n324_o & n327_o;
  /* HUC6280.vhd:296:24  */
  assign n329_o = n328_o ? 1'b1 : 1'b0;
  /* HUC6280.vhd:313:27  */
  assign n331_o = iop_sel | int_sel;
  /* HUC6280.vhd:313:38  */
  assign n332_o = n331_o | tmr_sel;
  /* HUC6280.vhd:313:49  */
  assign n333_o = n332_o | psg_sel;
  /* HUC6280.vhd:316:26  */
  assign n336_o = ~RST_N;
  /* HUC6280.vhd:321:53  */
  assign n338_o = ~cpu_we_n;
  /* HUC6280.vhd:321:41  */
  assign n339_o = n338_o ? cpu_do : cpu_di;
  /* HUC6280.vhd:319:25  */
  assign n341_o = en & io_sel;
  /* HUC6280.vhd:334:35  */
  assign n349_o = ~io_sel;
  /* HUC6280.vhd:341:43  */
  assign n350_o = cpu_a[1:0];
  /* HUC6280.vhd:343:65  */
  assign n351_o = io_buf[7:3];
  /* HUC6280.vhd:343:78  */
  assign n352_o = {n351_o, int_mask};
  /* HUC6280.vhd:342:41  */
  assign n354_o = n350_o == 2'b10;
  /* HUC6280.vhd:345:65  */
  assign n355_o = io_buf[7:3];
  /* HUC6280.vhd:345:78  */
  assign n356_o = {n355_o, tmr_irq};
  /* HUC6280.vhd:345:90  */
  assign n357_o = ~IRQ1_N;
  /* HUC6280.vhd:345:88  */
  assign n358_o = {n356_o, n357_o};
  /* HUC6280.vhd:345:103  */
  assign n359_o = ~IRQ2_N;
  /* HUC6280.vhd:345:101  */
  assign n360_o = {n358_o, n359_o};
  /* HUC6280.vhd:344:41  */
  assign n362_o = n350_o == 2'b11;
  assign n363_o = {n362_o, n354_o};
  /* HUC6280.vhd:341:33  */
  always @*
    case (n363_o)
      2'b10: n364_o = n360_o;
      2'b01: n364_o = n352_o;
      default: n364_o = io_buf;
    endcase
  /* HUC6280.vhd:350:49  */
  assign n365_o = io_buf[7];
  /* HUC6280.vhd:350:53  */
  assign n366_o = {n365_o, tmr_value};
  /* HUC6280.vhd:349:25  */
  assign n367_o = tmr_sel ? n366_o : io_buf;
  /* HUC6280.vhd:340:25  */
  assign n368_o = int_sel ? n364_o : n367_o;
  /* HUC6280.vhd:338:25  */
  assign n369_o = iop_sel ? K : n368_o;
  /* HUC6280.vhd:336:25  */
  assign n371_o = psg_sel ? 8'b00000000 : n369_o;
  /* HUC6280.vhd:334:25  */
  assign n372_o = n349_o ? DI : n371_o;
  /* HUC6280.vhd:97:17  */
  always @(posedge CLK or posedge n17_o)
    if (n17_o)
      n375_q <= 1'b0;
    else
      n375_q <= n46_o;
  /* HUC6280.vhd:97:17  */
  always @(posedge CLK or posedge n17_o)
    if (n17_o)
      n376_q <= 1'b0;
    else
      n376_q <= n53_o;
  /* HUC6280.vhd:97:17  */
  always @(posedge CLK or posedge n17_o)
    if (n17_o)
      n377_q <= 1'b0;
    else
      n377_q <= n61_o;
  /* HUC6280.vhd:333:17  */
  always @(posedge CLK)
    n378_q <= n372_o;
  /* HUC6280.vhd:167:17  */
  always @(posedge CLK or posedge n126_o)
    if (n126_o)
      n379_q <= 1'b1;
    else
      n379_q <= n146_o;
  /* HUC6280.vhd:97:17  */
  always @(posedge CLK or posedge n17_o)
    if (n17_o)
      n380_q <= 5'b00000;
    else
      n380_q <= n48_o;
  /* HUC6280.vhd:97:17  */
  always @(posedge CLK or posedge n17_o)
    if (n17_o)
      n381_q <= 3'b000;
    else
      n381_q <= n64_o;
  /* HUC6280.vhd:167:17  */
  assign n382_o = cpu_cer ? n131_o : vdc_sel_old;
  /* HUC6280.vhd:167:17  */
  always @(posedge CLK or posedge n126_o)
    if (n126_o)
      n383_q <= 1'b0;
    else
      n383_q <= n382_o;
  /* HUC6280.vhd:318:17  */
  assign n384_o = n341_o ? n339_o : io_buf;
  /* HUC6280.vhd:318:17  */
  always @(posedge CLK or posedge n336_o)
    if (n336_o)
      n385_q <= 8'b11111111;
    else
      n385_q <= n384_o;
  /* HUC6280.vhd:222:17  */
  assign n386_o = n226_o ? n214_o : int_mask;
  /* HUC6280.vhd:222:17  */
  always @(posedge CLK or posedge n203_o)
    if (n203_o)
      n387_q <= 3'b000;
    else
      n387_q <= n386_o;
  /* HUC6280.vhd:256:17  */
  always @(posedge CLK or posedge n249_o)
    if (n249_o)
      n388_q <= 10'b1111111111;
    else
      n388_q <= n291_o;
  /* HUC6280.vhd:256:17  */
  always @(posedge CLK or posedge n249_o)
    if (n249_o)
      n389_q <= 7'b0000000;
    else
      n389_q <= n299_o;
  /* HUC6280.vhd:256:17  */
  assign n390_o = n270_o ? n256_o : tmr_latch;
  /* HUC6280.vhd:256:17  */
  always @(posedge CLK or posedge n249_o)
    if (n249_o)
      n391_q <= 7'b0000000;
    else
      n391_q <= n390_o;
  /* HUC6280.vhd:256:17  */
  assign n392_o = n253_o ? n267_o : tmr_en;
  /* HUC6280.vhd:256:17  */
  always @(posedge CLK or posedge n249_o)
    if (n249_o)
      n393_q <= 1'b0;
    else
      n393_q <= n392_o;
  /* HUC6280.vhd:256:17  */
  assign n394_o = io_ce ? n294_o : tmr_reload;
  /* HUC6280.vhd:256:17  */
  always @(posedge CLK or posedge n249_o)
    if (n249_o)
      n395_q <= 1'b0;
    else
      n395_q <= n394_o;
  /* HUC6280.vhd:256:17  */
  always @(posedge CLK or posedge n249_o)
    if (n249_o)
      n396_q <= 1'b0;
    else
      n396_q <= n286_o;
  /* HUC6280.vhd:222:17  */
  always @(posedge CLK or posedge n203_o)
    if (n203_o)
      n397_q <= 1'b0;
    else
      n397_q <= n228_o;
  /* HUC6280.vhd:97:17  */
  always @(posedge CLK or posedge n17_o)
    if (n17_o)
      n398_q <= 1'b0;
    else
      n398_q <= n29_o;
  /* HUC6280.vhd:167:17  */
  always @(posedge CLK or posedge n126_o)
    if (n126_o)
      n399_q <= 1'b1;
    else
      n399_q <= n144_o;
  /* HUC6280.vhd:167:17  */
  always @(posedge CLK or posedge n126_o)
    if (n126_o)
      n400_q <= 1'b1;
    else
      n400_q <= n145_o;
  /* HUC6280.vhd:206:17  */
  assign n401_o = n186_o ? cpu_do : n402_q;
  /* HUC6280.vhd:206:17  */
  always @(posedge CLK or posedge n181_o)
    if (n181_o)
      n402_q <= 8'b00000000;
    else
      n402_q <= n401_o;
endmodule

