// common definitions used on tests
localparam TW=16;    // tone output bit width

// registers
localparam ATIME1=8,
           ATIME2=9,
           DTIME1=10,
           DTIME2=11,
           GCTL1 =12,
           GCTL2 =13;