module t48_int
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  [2:0] clk_mstate_i,
   input  jtf_executed_i,
   input  tim_overflow_i,
   input  en_tcnti_i,
   input  dis_tcnti_i,
   input  int_n_i,
   input  ale_i,
   input  last_cycle_i,
   input  en_i_i,
   input  dis_i_i,
   input  retr_executed_i,
   input  int_executed_i,
   output tf_o,
   output ext_int_o,
   output tim_int_o,
   output int_pending_o,
   output int_in_progress_o);
  wire [1:0] int_state_s;
  wire [1:0] int_state_q;
  wire timer_flag_q;
  wire timer_overflow_q;
  wire timer_int_enable_q;
  wire int_q;
  wire int_enable_q;
  wire ale_q;
  wire int_type_q;
  wire int_in_progress_q;
  wire n5070_o;
  wire n5072_o;
  wire n5073_o;
  wire [1:0] n5075_o;
  wire n5077_o;
  wire [1:0] n5079_o;
  wire n5081_o;
  wire [1:0] n5083_o;
  wire n5085_o;
  wire [2:0] n5086_o;
  reg [1:0] n5088_o;
  wire n5091_o;
  wire n5094_o;
  wire n5096_o;
  wire n5097_o;
  wire n5098_o;
  wire n5099_o;
  wire n5100_o;
  wire n5102_o;
  wire n5104_o;
  wire n5106_o;
  wire n5108_o;
  wire n5110_o;
  wire n5112_o;
  wire n5113_o;
  wire n5114_o;
  wire n5115_o;
  wire n5117_o;
  wire n5124_o;
  wire n5125_o;
  wire n5126_o;
  wire n5128_o;
  wire n5129_o;
  wire n5131_o;
  wire n5162_o;
  wire n5164_o;
  wire n5165_o;
  wire n5166_o;
  wire n5174_o;
  wire n5175_o;
  wire n5177_o;
  wire n5193_o;
  wire n5194_o;
  wire n5196_o;
  wire n5198_o;
  wire n5199_o;
  wire [1:0] n5200_o;
  reg [1:0] n5201_q;
  wire n5202_o;
  reg n5203_q;
  wire n5204_o;
  reg n5205_q;
  wire n5206_o;
  reg n5207_q;
  wire n5208_o;
  reg n5209_q;
  wire n5210_o;
  reg n5211_q;
  wire n5212_o;
  reg n5213_q;
  wire n5214_o;
  reg n5215_q;
  wire n5216_o;
  reg n5217_q;
  assign tf_o = n5193_o;
  assign ext_int_o = int_type_q;
  assign tim_int_o = n5194_o;
  assign int_pending_o = n5196_o;
  assign int_in_progress_o = n5199_o;
  /* int.vhd:91:10  */
  assign int_state_s = n5088_o; // (signal)
  /* int.vhd:92:10  */
  assign int_state_q = n5201_q; // (signal)
  /* int.vhd:94:10  */
  assign timer_flag_q = n5203_q; // (signal)
  /* int.vhd:95:10  */
  assign timer_overflow_q = n5205_q; // (signal)
  /* int.vhd:96:10  */
  assign timer_int_enable_q = n5207_q; // (signal)
  /* int.vhd:97:10  */
  assign int_q = n5209_q; // (signal)
  /* int.vhd:98:10  */
  assign int_enable_q = n5211_q; // (signal)
  /* int.vhd:99:10  */
  assign ale_q = n5213_q; // (signal)
  /* int.vhd:100:10  */
  assign int_type_q = n5215_q; // (signal)
  /* int.vhd:101:10  */
  assign int_in_progress_q = n5217_q; // (signal)
  /* int.vhd:123:30  */
  assign n5070_o = int_in_progress_q & last_cycle_i;
  /* int.vhd:124:42  */
  assign n5072_o = clk_mstate_i == 3'b100;
  /* int.vhd:124:25  */
  assign n5073_o = n5070_o & n5072_o;
  /* int.vhd:123:9  */
  assign n5075_o = n5073_o ? 2'b01 : int_state_q;
  /* int.vhd:122:7  */
  assign n5077_o = int_state_q == 2'b00;
  /* int.vhd:129:9  */
  assign n5079_o = int_executed_i ? 2'b10 : int_state_q;
  /* int.vhd:128:7  */
  assign n5081_o = int_state_q == 2'b01;
  /* int.vhd:134:9  */
  assign n5083_o = retr_executed_i ? 2'b00 : int_state_q;
  /* int.vhd:133:7  */
  assign n5085_o = int_state_q == 2'b10;
  assign n5086_o = {n5085_o, n5081_o, n5077_o};
  /* int.vhd:121:5  */
  always @*
    case (n5086_o)
      3'b100: n5088_o = n5083_o;
      3'b010: n5088_o = n5079_o;
      3'b001: n5088_o = n5075_o;
      default: n5088_o = 2'b00;
    endcase
  /* int.vhd:158:14  */
  assign n5091_o = ~res_i;
  /* int.vhd:174:9  */
  assign n5094_o = tim_overflow_i ? 1'b1 : timer_flag_q;
  /* int.vhd:172:9  */
  assign n5096_o = jtf_executed_i ? 1'b0 : n5094_o;
  /* int.vhd:178:24  */
  assign n5097_o = ~int_type_q;
  /* int.vhd:178:36  */
  assign n5098_o = n5097_o & int_executed_i;
  /* int.vhd:179:11  */
  assign n5099_o = ~timer_int_enable_q;
  /* int.vhd:178:56  */
  assign n5100_o = n5098_o | n5099_o;
  /* int.vhd:181:9  */
  assign n5102_o = tim_overflow_i ? 1'b1 : timer_overflow_q;
  /* int.vhd:178:9  */
  assign n5104_o = n5100_o ? 1'b0 : n5102_o;
  /* int.vhd:187:9  */
  assign n5106_o = en_tcnti_i ? 1'b1 : timer_int_enable_q;
  /* int.vhd:185:9  */
  assign n5108_o = dis_tcnti_i ? 1'b0 : n5106_o;
  /* int.vhd:193:9  */
  assign n5110_o = en_i_i ? 1'b1 : int_enable_q;
  /* int.vhd:191:9  */
  assign n5112_o = dis_i_i ? 1'b0 : n5110_o;
  /* int.vhd:199:22  */
  assign n5113_o = int_q & int_enable_q;
  /* int.vhd:199:40  */
  assign n5114_o = n5113_o | timer_overflow_q;
  /* int.vhd:202:14  */
  assign n5115_o = ~int_in_progress_q;
  /* int.vhd:203:45  */
  assign n5117_o = int_q & int_enable_q;
  /* t48_pack-p.vhd:66:5  */
  assign n5124_o = n5117_o ? 1'b1 : 1'b0;
  /* int.vhd:199:9  */
  assign n5125_o = n5126_o ? n5124_o : int_type_q;
  /* int.vhd:199:9  */
  assign n5126_o = n5114_o & n5115_o;
  /* int.vhd:199:9  */
  assign n5128_o = n5114_o ? 1'b1 : int_in_progress_q;
  /* int.vhd:197:9  */
  assign n5129_o = retr_executed_i ? int_type_q : n5125_o;
  /* int.vhd:197:9  */
  assign n5131_o = retr_executed_i ? 1'b0 : n5128_o;
  /* int.vhd:224:14  */
  assign n5162_o = ~res_i;
  /* int.vhd:232:25  */
  assign n5164_o = last_cycle_i & ale_q;
  /* int.vhd:233:22  */
  assign n5165_o = ~ale_i;
  /* int.vhd:233:18  */
  assign n5166_o = n5164_o & n5165_o;
  /* t48_pack-p.vhd:75:5  */
  assign n5174_o = int_n_i ? 1'b1 : 1'b0;
  /* int.vhd:234:20  */
  assign n5175_o = ~n5174_o;
  /* int.vhd:229:7  */
  assign n5177_o = xtal_en_i & n5166_o;
  /* t48_pack-p.vhd:66:5  */
  assign n5193_o = timer_flag_q ? 1'b1 : 1'b0;
  /* int.vhd:249:35  */
  assign n5194_o = ~int_type_q;
  /* int.vhd:250:36  */
  assign n5196_o = int_state_q == 2'b01;
  /* int.vhd:251:58  */
  assign n5198_o = int_state_q != 2'b00;
  /* int.vhd:251:42  */
  assign n5199_o = int_in_progress_q & n5198_o;
  /* int.vhd:167:5  */
  assign n5200_o = en_clk_i ? int_state_s : int_state_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n5091_o)
    if (n5091_o)
      n5201_q <= 2'b00;
    else
      n5201_q <= n5200_o;
  /* int.vhd:167:5  */
  assign n5202_o = en_clk_i ? n5096_o : timer_flag_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n5091_o)
    if (n5091_o)
      n5203_q <= 1'b0;
    else
      n5203_q <= n5202_o;
  /* int.vhd:167:5  */
  assign n5204_o = en_clk_i ? n5104_o : timer_overflow_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n5091_o)
    if (n5091_o)
      n5205_q <= 1'b0;
    else
      n5205_q <= n5204_o;
  /* int.vhd:167:5  */
  assign n5206_o = en_clk_i ? n5108_o : timer_int_enable_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n5091_o)
    if (n5091_o)
      n5207_q <= 1'b0;
    else
      n5207_q <= n5206_o;
  /* int.vhd:228:5  */
  assign n5208_o = n5177_o ? n5175_o : int_q;
  /* int.vhd:228:5  */
  always @(posedge xtal_i or posedge n5162_o)
    if (n5162_o)
      n5209_q <= 1'b0;
    else
      n5209_q <= n5208_o;
  /* int.vhd:167:5  */
  assign n5210_o = en_clk_i ? n5112_o : int_enable_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n5091_o)
    if (n5091_o)
      n5211_q <= 1'b0;
    else
      n5211_q <= n5210_o;
  /* int.vhd:228:5  */
  assign n5212_o = xtal_en_i ? ale_i : ale_q;
  /* int.vhd:228:5  */
  always @(posedge xtal_i or posedge n5162_o)
    if (n5162_o)
      n5213_q <= 1'b0;
    else
      n5213_q <= n5212_o;
  /* int.vhd:167:5  */
  assign n5214_o = en_clk_i ? n5129_o : int_type_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n5091_o)
    if (n5091_o)
      n5215_q <= 1'b0;
    else
      n5215_q <= n5214_o;
  /* int.vhd:167:5  */
  assign n5216_o = en_clk_i ? n5131_o : int_in_progress_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n5091_o)
    if (n5091_o)
      n5217_q <= 1'b0;
    else
      n5217_q <= n5216_o;
endmodule

module t48_psw
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  read_psw_i,
   input  read_sp_i,
   input  write_psw_i,
   input  write_sp_i,
   input  special_data_i,
   input  inc_stackp_i,
   input  dec_stackp_i,
   input  write_carry_i,
   input  write_aux_carry_i,
   input  write_f0_i,
   input  write_bs_i,
   input  aux_carry_i,
   output [7:0] data_o,
   output carry_o,
   output aux_carry_o,
   output f0_o,
   output bs_o);
  wire [3:0] psw_q;
  wire [2:0] sp_q;
  wire n5002_o;
  wire [2:0] n5006_o;
  wire [2:0] n5007_o;
  wire [2:0] n5009_o;
  wire [2:0] n5010_o;
  wire [2:0] n5012_o;
  wire [2:0] n5013_o;
  wire n5014_o;
  wire n5015_o;
  wire n5016_o;
  wire n5017_o;
  wire n5021_o;
  wire n5022_o;
  wire n5023_o;
  wire n5024_o;
  wire n5028_o;
  wire n5029_o;
  wire n5030_o;
  wire n5031_o;
  wire n5032_o;
  wire n5033_o;
  wire n5034_o;
  wire n5035_o;
  wire [3:0] n5036_o;
  wire [3:0] n5048_o;
  localparam [7:0] n5049_o = 8'b11111111;
  wire [3:0] n5050_o;
  wire [3:0] n5052_o;
  wire [3:0] n5053_o;
  wire n5055_o;
  wire n5056_o;
  wire n5057_o;
  wire n5058_o;
  wire [3:0] n5059_o;
  reg [3:0] n5060_q;
  wire [2:0] n5061_o;
  reg [2:0] n5062_q;
  wire [7:0] n5063_o;
  assign data_o = n5063_o;
  assign carry_o = n5055_o;
  assign aux_carry_o = n5056_o;
  assign f0_o = n5057_o;
  assign bs_o = n5058_o;
  /* psw.vhd:101:10  */
  assign psw_q = n5060_q; // (signal)
  /* psw.vhd:103:10  */
  assign sp_q = n5062_q; // (signal)
  /* psw.vhd:119:14  */
  assign n5002_o = ~res_i;
  /* psw.vhd:131:34  */
  assign n5006_o = data_i[2:0];
  /* psw.vhd:130:9  */
  assign n5007_o = write_sp_i ? n5006_o : sp_q;
  /* psw.vhd:136:25  */
  assign n5009_o = sp_q + 3'b001;
  /* psw.vhd:135:9  */
  assign n5010_o = inc_stackp_i ? n5009_o : n5007_o;
  /* psw.vhd:140:25  */
  assign n5012_o = sp_q - 3'b001;
  /* psw.vhd:139:9  */
  assign n5013_o = dec_stackp_i ? n5012_o : n5010_o;
  assign n5014_o = data_i[7];
  assign n5015_o = psw_q[3];
  /* psw.vhd:127:9  */
  assign n5016_o = write_psw_i ? n5014_o : n5015_o;
  /* psw.vhd:144:9  */
  assign n5017_o = write_carry_i ? special_data_i : n5016_o;
  assign n5021_o = data_i[6];
  assign n5022_o = psw_q[2];
  /* psw.vhd:127:9  */
  assign n5023_o = write_psw_i ? n5021_o : n5022_o;
  /* psw.vhd:148:9  */
  assign n5024_o = write_aux_carry_i ? aux_carry_i : n5023_o;
  assign n5028_o = data_i[5];
  assign n5029_o = psw_q[1];
  /* psw.vhd:127:9  */
  assign n5030_o = write_psw_i ? n5028_o : n5029_o;
  /* psw.vhd:152:9  */
  assign n5031_o = write_f0_i ? special_data_i : n5030_o;
  assign n5032_o = data_i[4];
  assign n5033_o = psw_q[0];
  /* psw.vhd:127:9  */
  assign n5034_o = write_psw_i ? n5032_o : n5033_o;
  /* psw.vhd:156:9  */
  assign n5035_o = write_bs_i ? special_data_i : n5034_o;
  assign n5036_o = {n5017_o, n5024_o, n5031_o, n5035_o};
  /* psw.vhd:182:5  */
  assign n5048_o = read_psw_i ? psw_q : 4'b1111;
  assign n5050_o = n5049_o[3:0];
  /* psw.vhd:187:33  */
  assign n5052_o = {1'b1, sp_q};
  /* psw.vhd:186:5  */
  assign n5053_o = read_sp_i ? n5052_o : n5050_o;
  /* psw.vhd:207:23  */
  assign n5055_o = psw_q[3];
  /* psw.vhd:208:23  */
  assign n5056_o = psw_q[2];
  /* psw.vhd:209:23  */
  assign n5057_o = psw_q[1];
  /* psw.vhd:210:23  */
  assign n5058_o = psw_q[0];
  /* psw.vhd:123:5  */
  assign n5059_o = en_clk_i ? n5036_o : psw_q;
  /* psw.vhd:123:5  */
  always @(posedge clk_i or posedge n5002_o)
    if (n5002_o)
      n5060_q <= 4'b0000;
    else
      n5060_q <= n5059_o;
  /* psw.vhd:123:5  */
  assign n5061_o = en_clk_i ? n5013_o : sp_q;
  /* psw.vhd:123:5  */
  always @(posedge clk_i or posedge n5002_o)
    if (n5002_o)
      n5062_q <= 3'b000;
    else
      n5062_q <= n5061_o;
  /* psw.vhd:119:5  */
  assign n5063_o = {n5048_o, n5053_o};
endmodule

module t48_pmem_ctrl
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_pcl_i,
   input  read_pcl_i,
   input  write_pch_i,
   input  read_pch_i,
   input  inc_pc_i,
   input  write_pmem_addr_i,
   input  [1:0] addr_type_i,
   input  read_pmem_i,
   input  [7:0] pmem_data_i,
   output [7:0] data_o,
   output [11:0] pmem_addr_o);
  wire [11:0] program_counter_q;
  wire [11:0] pmem_addr_s;
  wire [11:0] pmem_addr_q;
  wire n4928_o;
  wire [3:0] n4930_o;
  wire [10:0] n4931_o;
  wire [10:0] n4933_o;
  wire [10:0] n4934_o;
  wire [10:0] n4935_o;
  wire [7:0] n4936_o;
  wire [7:0] n4937_o;
  wire [7:0] n4938_o;
  wire [2:0] n4939_o;
  wire [2:0] n4940_o;
  wire [2:0] n4941_o;
  wire n4942_o;
  wire n4943_o;
  wire n4944_o;
  wire [11:0] n4945_o;
  wire [7:0] n4946_o;
  wire [7:0] n4947_o;
  wire [3:0] n4948_o;
  wire [3:0] n4949_o;
  wire [3:0] n4950_o;
  wire [11:0] n4952_o;
  wire n4954_o;
  wire n4964_o;
  wire n4966_o;
  wire n4969_o;
  wire [2:0] n4970_o;
  wire [7:0] n4971_o;
  reg [7:0] n4972_o;
  wire [3:0] n4973_o;
  reg [3:0] n4974_o;
  wire [7:0] n4978_o;
  wire [3:0] n4979_o;
  wire [3:0] n4981_o;
  wire [3:0] n4982_o;
  wire [3:0] n4983_o;
  wire [3:0] n4984_o;
  wire [3:0] n4986_o;
  wire [7:0] n4987_o;
  wire [7:0] n4988_o;
  wire [11:0] n4991_o;
  reg [11:0] n4992_q;
  wire [11:0] n4993_o;
  wire [11:0] n4994_o;
  reg [11:0] n4995_q;
  assign data_o = n4988_o;
  assign pmem_addr_o = pmem_addr_q;
  /* pmem_ctrl.vhd:98:10  */
  assign program_counter_q = n4992_q; // (signal)
  /* pmem_ctrl.vhd:102:10  */
  assign pmem_addr_s = n4993_o; // (signal)
  /* pmem_ctrl.vhd:103:10  */
  assign pmem_addr_q = n4995_q; // (signal)
  /* pmem_ctrl.vhd:115:14  */
  assign n4928_o = ~res_i;
  /* pmem_ctrl.vhd:127:28  */
  assign n4930_o = data_i[3:0];
  /* pmem_ctrl.vhd:133:30  */
  assign n4931_o = program_counter_q[10:0];
  /* pmem_ctrl.vhd:133:49  */
  assign n4933_o = n4931_o + 11'b00000000001;
  /* p2.vhd:153:3  */
  assign n4934_o = program_counter_q[10:0];
  /* pmem_ctrl.vhd:128:9  */
  assign n4935_o = inc_pc_i ? n4933_o : n4934_o;
  /* p2.vhd:115:5  */
  assign n4936_o = n4935_o[7:0];
  /* p2.vhd:115:5  */
  assign n4937_o = program_counter_q[7:0];
  /* pmem_ctrl.vhd:125:9  */
  assign n4938_o = write_pch_i ? n4937_o : n4936_o;
  /* decoder.vhd:521:15  */
  assign n4939_o = n4935_o[10:8];
  /* decoder.vhd:521:15  */
  assign n4940_o = n4930_o[2:0];
  /* pmem_ctrl.vhd:125:9  */
  assign n4941_o = write_pch_i ? n4940_o : n4939_o;
  /* p2.vhd:155:5  */
  assign n4942_o = n4930_o[3];
  assign n4943_o = program_counter_q[11];
  /* pmem_ctrl.vhd:125:9  */
  assign n4944_o = write_pch_i ? n4942_o : n4943_o;
  /* decoder_pack-p.vhd:116:14  */
  assign n4945_o = {n4944_o, n4941_o, n4938_o};
  assign n4946_o = n4945_o[7:0];
  /* pmem_ctrl.vhd:123:9  */
  assign n4947_o = write_pcl_i ? data_i : n4946_o;
  assign n4948_o = n4945_o[11:8];
  /* decoder_pack-p.vhd:114:14  */
  assign n4949_o = program_counter_q[11:8];
  /* pmem_ctrl.vhd:123:9  */
  assign n4950_o = write_pcl_i ? n4949_o : n4948_o;
  /* decoder_pack-p.vhd:112:12  */
  assign n4952_o = {n4950_o, n4947_o};
  /* pmem_ctrl.vhd:120:7  */
  assign n4954_o = en_clk_i & write_pmem_addr_i;
  /* pmem_ctrl.vhd:165:7  */
  assign n4964_o = addr_type_i == 2'b00;
  /* pmem_ctrl.vhd:169:7  */
  assign n4966_o = addr_type_i == 2'b01;
  /* pmem_ctrl.vhd:175:7  */
  assign n4969_o = addr_type_i == 2'b10;
  /* decoder_pack-p.vhd:545:14  */
  assign n4970_o = {n4969_o, n4966_o, n4964_o};
  assign n4971_o = program_counter_q[7:0];
  /* pmem_ctrl.vhd:164:5  */
  always @*
    case (n4970_o)
      3'b100: n4972_o = data_i;
      3'b010: n4972_o = data_i;
      3'b001: n4972_o = n4971_o;
      default: n4972_o = n4971_o;
    endcase
  assign n4973_o = program_counter_q[11:8];
  /* pmem_ctrl.vhd:164:5  */
  always @*
    case (n4970_o)
      3'b100: n4974_o = 4'b0011;
      3'b010: n4974_o = n4973_o;
      3'b001: n4974_o = n4973_o;
      default: n4974_o = n4973_o;
    endcase
  /* pmem_ctrl.vhd:207:51  */
  assign n4978_o = program_counter_q[7:0];
  /* pmem_ctrl.vhd:209:63  */
  assign n4979_o = program_counter_q[11:8];
  /* pmem_ctrl.vhd:208:5  */
  assign n4981_o = read_pch_i ? n4979_o : 4'b1111;
  assign n4982_o = n4978_o[3:0];
  /* pmem_ctrl.vhd:206:5  */
  assign n4983_o = read_pcl_i ? n4982_o : n4981_o;
  assign n4984_o = n4978_o[7:4];
  /* pmem_ctrl.vhd:206:5  */
  assign n4986_o = read_pcl_i ? n4984_o : 4'b1111;
  assign n4987_o = {n4986_o, n4983_o};
  /* pmem_ctrl.vhd:204:5  */
  assign n4988_o = read_pmem_i ? pmem_data_i : n4987_o;
  /* pmem_ctrl.vhd:119:5  */
  assign n4991_o = en_clk_i ? n4952_o : program_counter_q;
  /* pmem_ctrl.vhd:119:5  */
  always @(posedge clk_i or posedge n4928_o)
    if (n4928_o)
      n4992_q <= 12'b000000000000;
    else
      n4992_q <= n4991_o;
  /* pmem_ctrl.vhd:115:5  */
  assign n4993_o = {n4974_o, n4972_o};
  /* pmem_ctrl.vhd:119:5  */
  assign n4994_o = n4954_o ? pmem_addr_s : pmem_addr_q;
  /* pmem_ctrl.vhd:119:5  */
  always @(posedge clk_i or posedge n4928_o)
    if (n4928_o)
      n4995_q <= 12'b000000000000;
    else
      n4995_q <= n4994_o;
endmodule

module t48_p2
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  [7:0] data_i,
   input  write_p2_i,
   input  write_exp_i,
   input  read_p2_i,
   input  read_reg_i,
   input  read_exp_i,
   input  output_pch_i,
   input  [3:0] pch_i,
   input  [7:0] p2_i,
   output [7:0] data_o,
   output [7:0] p2_o,
   output p2l_low_imp_o,
   output p2h_low_imp_o);
  wire [7:0] p2_q;
  wire l_low_imp_q;
  wire h_low_imp_q;
  wire en_clk_q;
  wire l_low_imp_del_q;
  wire h_low_imp_del_q;
  wire output_pch_q;
  wire n4827_o;
  wire [3:0] n4829_o;
  wire [3:0] n4830_o;
  wire [3:0] n4831_o;
  wire n4834_o;
  wire [3:0] n4835_o;
  wire [3:0] n4836_o;
  wire [3:0] n4837_o;
  wire [3:0] n4838_o;
  wire [3:0] n4839_o;
  wire n4841_o;
  wire n4845_o;
  wire [7:0] n4847_o;
  wire n4862_o;
  wire [3:0] n4864_o;
  wire [3:0] n4865_o;
  wire [3:0] n4866_o;
  wire n4867_o;
  wire n4868_o;
  wire n4869_o;
  wire n4872_o;
  wire n4873_o;
  wire n4876_o;
  wire [7:0] n4877_o;
  wire [3:0] n4900_o;
  wire [7:0] n4902_o;
  wire [7:0] n4903_o;
  wire [7:0] n4904_o;
  wire [7:0] n4906_o;
  wire [7:0] n4909_o;
  reg [7:0] n4910_q;
  wire n4911_o;
  reg n4912_q;
  wire n4913_o;
  reg n4914_q;
  wire n4915_o;
  reg n4916_q;
  wire n4917_o;
  reg n4918_q;
  wire n4919_o;
  reg n4920_q;
  wire n4921_o;
  reg n4922_q;
  wire [7:0] n4923_o;
  reg [7:0] n4924_q;
  assign data_o = n4906_o;
  assign p2_o = n4924_q;
  assign p2l_low_imp_o = l_low_imp_del_q;
  assign p2h_low_imp_o = h_low_imp_del_q;
  /* p2.vhd:89:10  */
  assign p2_q = n4910_q; // (signal)
  /* p2.vhd:92:10  */
  assign l_low_imp_q = n4912_q; // (signal)
  /* p2.vhd:93:10  */
  assign h_low_imp_q = n4914_q; // (signal)
  /* p2.vhd:95:10  */
  assign en_clk_q = n4916_q; // (signal)
  /* p2.vhd:96:10  */
  assign l_low_imp_del_q = n4918_q; // (signal)
  /* p2.vhd:97:10  */
  assign h_low_imp_del_q = n4920_q; // (signal)
  /* p2.vhd:98:10  */
  assign output_pch_q = n4922_q; // (signal)
  /* p2.vhd:110:14  */
  assign n4827_o = ~res_i;
  /* p2.vhd:129:41  */
  assign n4829_o = data_i[3:0];
  /* decoder.vhd:496:15  */
  assign n4830_o = p2_q[3:0];
  /* p2.vhd:127:9  */
  assign n4831_o = write_exp_i ? n4829_o : n4830_o;
  /* p2.vhd:127:9  */
  assign n4834_o = write_exp_i ? 1'b1 : 1'b0;
  /* decoder.vhd:521:15  */
  assign n4835_o = data_i[3:0];
  /* p2.vhd:121:9  */
  assign n4836_o = write_p2_i ? n4835_o : n4831_o;
  /* decoder.vhd:521:15  */
  assign n4837_o = data_i[7:4];
  /* decoder.vhd:521:15  */
  assign n4838_o = p2_q[7:4];
  /* p2.vhd:121:9  */
  assign n4839_o = write_p2_i ? n4837_o : n4838_o;
  /* p2.vhd:121:9  */
  assign n4841_o = write_p2_i ? 1'b1 : n4834_o;
  /* p2.vhd:121:9  */
  assign n4845_o = write_p2_i ? 1'b1 : 1'b0;
  assign n4847_o = {n4839_o, n4836_o};
  /* p2.vhd:155:14  */
  assign n4862_o = ~res_i;
  /* decoder.vhd:506:15  */
  assign n4864_o = p2_q[3:0];
  /* p2.vhd:170:9  */
  assign n4865_o = output_pch_i ? pch_i : n4864_o;
  /* decoder.vhd:499:26  */
  assign n4866_o = p2_q[7:4];
  /* p2.vhd:179:26  */
  assign n4867_o = output_pch_q ^ output_pch_i;
  /* p2.vhd:179:44  */
  assign n4868_o = n4867_o | l_low_imp_q;
  /* p2.vhd:178:21  */
  assign n4869_o = en_clk_q & n4868_o;
  /* p2.vhd:178:9  */
  assign n4872_o = n4869_o ? 1'b1 : 1'b0;
  /* p2.vhd:189:21  */
  assign n4873_o = en_clk_q & h_low_imp_q;
  /* p2.vhd:189:9  */
  assign n4876_o = n4873_o ? 1'b1 : 1'b0;
  /* decoder.vhd:499:22  */
  assign n4877_o = {n4866_o, n4865_o};
  /* p2.vhd:221:32  */
  assign n4900_o = p2_i[3:0];
  /* p2.vhd:221:26  */
  assign n4902_o = {4'b0000, n4900_o};
  /* p2.vhd:220:7  */
  assign n4903_o = read_exp_i ? n4902_o : p2_i;
  /* p2.vhd:218:7  */
  assign n4904_o = read_reg_i ? p2_q : n4903_o;
  /* p2.vhd:217:5  */
  assign n4906_o = read_p2_i ? n4904_o : 8'b11111111;
  /* p2.vhd:115:5  */
  assign n4909_o = en_clk_i ? n4847_o : p2_q;
  /* p2.vhd:115:5  */
  always @(posedge clk_i or posedge n4827_o)
    if (n4827_o)
      n4910_q <= 8'b11111111;
    else
      n4910_q <= n4909_o;
  /* p2.vhd:115:5  */
  assign n4911_o = en_clk_i ? n4841_o : l_low_imp_q;
  /* p2.vhd:115:5  */
  always @(posedge clk_i or posedge n4827_o)
    if (n4827_o)
      n4912_q <= 1'b0;
    else
      n4912_q <= n4911_o;
  /* p2.vhd:115:5  */
  assign n4913_o = en_clk_i ? n4845_o : h_low_imp_q;
  /* p2.vhd:115:5  */
  always @(posedge clk_i or posedge n4827_o)
    if (n4827_o)
      n4914_q <= 1'b0;
    else
      n4914_q <= n4913_o;
  /* p2.vhd:162:5  */
  assign n4915_o = xtal_en_i ? en_clk_i : en_clk_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4862_o)
    if (n4862_o)
      n4916_q <= 1'b0;
    else
      n4916_q <= n4915_o;
  /* p2.vhd:162:5  */
  assign n4917_o = xtal_en_i ? n4872_o : l_low_imp_del_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4862_o)
    if (n4862_o)
      n4918_q <= 1'b0;
    else
      n4918_q <= n4917_o;
  /* p2.vhd:162:5  */
  assign n4919_o = xtal_en_i ? n4876_o : h_low_imp_del_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4862_o)
    if (n4862_o)
      n4920_q <= 1'b0;
    else
      n4920_q <= n4919_o;
  /* p2.vhd:162:5  */
  assign n4921_o = xtal_en_i ? output_pch_i : output_pch_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4862_o)
    if (n4862_o)
      n4922_q <= 1'b0;
    else
      n4922_q <= n4921_o;
  /* p2.vhd:162:5  */
  assign n4923_o = xtal_en_i ? n4877_o : n4924_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4862_o)
    if (n4862_o)
      n4924_q <= 8'b11111111;
    else
      n4924_q <= n4923_o;
endmodule

module t48_p1
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_p1_i,
   input  read_p1_i,
   input  read_reg_i,
   input  [7:0] p1_i,
   output [7:0] data_o,
   output [7:0] p1_o,
   output p1_low_imp_o);
  wire [7:0] p1_q;
  wire low_imp_q;
  wire n4797_o;
  wire n4802_o;
  wire n4803_o;
  wire [7:0] n4813_o;
  wire [7:0] n4815_o;
  wire [7:0] n4818_o;
  reg [7:0] n4819_q;
  wire n4820_o;
  reg n4821_q;
  assign data_o = n4815_o;
  assign p1_o = p1_q;
  assign p1_low_imp_o = low_imp_q;
  /* p1.vhd:81:10  */
  assign p1_q = n4819_q; // (signal)
  /* p1.vhd:84:10  */
  assign low_imp_q = n4821_q; // (signal)
  /* p1.vhd:96:14  */
  assign n4797_o = ~res_i;
  /* p1.vhd:103:9  */
  assign n4802_o = write_p1_i ? 1'b1 : 1'b0;
  /* p1.vhd:101:7  */
  assign n4803_o = en_clk_i & write_p1_i;
  /* p1.vhd:133:7  */
  assign n4813_o = read_reg_i ? p1_q : p1_i;
  /* p1.vhd:132:5  */
  assign n4815_o = read_p1_i ? n4813_o : 8'b11111111;
  /* p1.vhd:100:5  */
  assign n4818_o = n4803_o ? data_i : p1_q;
  /* p1.vhd:100:5  */
  always @(posedge clk_i or posedge n4797_o)
    if (n4797_o)
      n4819_q <= 8'b11111111;
    else
      n4819_q <= n4818_o;
  /* p1.vhd:100:5  */
  assign n4820_o = en_clk_i ? n4802_o : low_imp_q;
  /* p1.vhd:100:5  */
  always @(posedge clk_i or posedge n4797_o)
    if (n4797_o)
      n4821_q <= 1'b0;
    else
      n4821_q <= n4820_o;
endmodule

module t48_timer_4
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  t1_i,
   input  [2:0] clk_mstate_i,
   input  [7:0] data_i,
   input  read_timer_i,
   input  write_timer_i,
   input  start_t_i,
   input  start_cnt_i,
   input  stop_tcnt_i,
   output [7:0] data_o,
   output overflow_o);
  wire [7:0] counter_q;
  wire overflow_q;
  wire increment_s;
  wire [1:0] inc_sel_q;
  wire t1_q;
  wire t1_inc_s;
  wire [4:0] prescaler_q;
  wire pre_inc_s;
  wire n4683_o;
  wire n4685_o;
  wire n4687_o;
  wire n4688_o;
  wire n4689_o;
  wire n4692_o;
  wire n4694_o;
  wire n4698_o;
  wire n4700_o;
  wire n4701_o;
  wire n4704_o;
  wire n4706_o;
  wire n4708_o;
  wire [2:0] n4709_o;
  reg n4712_o;
  wire n4716_o;
  wire [7:0] n4719_o;
  wire n4721_o;
  wire n4724_o;
  wire [7:0] n4725_o;
  wire n4727_o;
  wire [7:0] n4728_o;
  wire n4730_o;
  wire n4733_o;
  wire n4735_o;
  wire n4737_o;
  wire n4740_o;
  wire [4:0] n4742_o;
  wire [4:0] n4743_o;
  wire [4:0] n4745_o;
  wire [1:0] n4747_o;
  wire [1:0] n4749_o;
  wire [1:0] n4751_o;
  wire n4755_o;
  wire [7:0] n4773_o;
  wire n4782_o;
  wire [7:0] n4783_o;
  reg [7:0] n4784_q;
  wire n4785_o;
  reg n4786_q;
  wire [1:0] n4787_o;
  reg [1:0] n4788_q;
  wire n4789_o;
  reg n4790_q;
  wire [4:0] n4791_o;
  reg [4:0] n4792_q;
  assign data_o = n4773_o;
  assign overflow_o = n4782_o;
  /* timer.vhd:89:10  */
  assign counter_q = n4784_q; // (signal)
  /* timer.vhd:90:10  */
  assign overflow_q = n4786_q; // (signal)
  /* timer.vhd:94:10  */
  assign increment_s = n4712_o; // (signal)
  /* timer.vhd:95:10  */
  assign inc_sel_q = n4788_q; // (signal)
  /* timer.vhd:98:10  */
  assign t1_q = n4790_q; // (signal)
  /* timer.vhd:99:10  */
  assign t1_inc_s = n4694_o; // (signal)
  /* timer.vhd:102:10  */
  assign prescaler_q = n4792_q; // (signal)
  /* timer.vhd:103:10  */
  assign pre_inc_s = n4701_o; // (signal)
  /* timer.vhd:134:48  */
  assign n4683_o = clk_mstate_i == 3'b011;
  /* timer.vhd:134:31  */
  assign n4685_o = 1'b1 & n4683_o;
  /* timer.vhd:133:59  */
  assign n4687_o = 1'b0 | n4685_o;
  /* timer.vhd:136:30  */
  assign n4688_o = ~t1_i;
  /* timer.vhd:136:21  */
  assign n4689_o = t1_q & n4688_o;
  /* timer.vhd:136:7  */
  assign n4692_o = n4689_o ? 1'b1 : 1'b0;
  /* timer.vhd:133:5  */
  assign n4694_o = n4687_o ? n4692_o : 1'b0;
  /* timer.vhd:146:29  */
  assign n4698_o = clk_mstate_i == 3'b011;
  /* timer.vhd:146:55  */
  assign n4700_o = prescaler_q == 5'b11111;
  /* timer.vhd:146:39  */
  assign n4701_o = n4698_o & n4700_o;
  /* timer.vhd:163:7  */
  assign n4704_o = inc_sel_q == 2'b00;
  /* timer.vhd:165:7  */
  assign n4706_o = inc_sel_q == 2'b01;
  /* timer.vhd:167:7  */
  assign n4708_o = inc_sel_q == 2'b10;
  assign n4709_o = {n4708_o, n4706_o, n4704_o};
  /* timer.vhd:162:5  */
  always @*
    case (n4709_o)
      3'b100: n4712_o = t1_inc_s;
      3'b010: n4712_o = pre_inc_s;
      3'b001: n4712_o = 1'b0;
      default: n4712_o = 1'b0;
    endcase
  /* timer.vhd:186:14  */
  assign n4716_o = ~res_i;
  /* timer.vhd:203:37  */
  assign n4719_o = counter_q + 8'b00000001;
  /* timer.vhd:205:24  */
  assign n4721_o = counter_q == 8'b11111111;
  /* timer.vhd:205:11  */
  assign n4724_o = n4721_o ? 1'b1 : 1'b0;
  /* timer.vhd:202:9  */
  assign n4725_o = increment_s ? n4719_o : counter_q;
  /* timer.vhd:202:9  */
  assign n4727_o = increment_s ? n4724_o : 1'b0;
  /* timer.vhd:199:9  */
  assign n4728_o = write_timer_i ? data_i : n4725_o;
  /* timer.vhd:199:9  */
  assign n4730_o = write_timer_i ? 1'b0 : n4727_o;
  /* timer.vhd:213:52  */
  assign n4733_o = clk_mstate_i == 3'b011;
  /* timer.vhd:213:35  */
  assign n4735_o = 1'b1 & n4733_o;
  /* timer.vhd:212:63  */
  assign n4737_o = 1'b0 | n4735_o;
  /* timer.vhd:221:28  */
  assign n4740_o = clk_mstate_i == 3'b010;
  /* timer.vhd:222:39  */
  assign n4742_o = prescaler_q + 5'b00001;
  /* timer.vhd:221:9  */
  assign n4743_o = n4740_o ? n4742_o : prescaler_q;
  /* timer.vhd:218:9  */
  assign n4745_o = start_t_i ? 5'b00000 : n4743_o;
  /* timer.vhd:231:9  */
  assign n4747_o = stop_tcnt_i ? 2'b00 : inc_sel_q;
  /* timer.vhd:229:9  */
  assign n4749_o = start_cnt_i ? 2'b10 : n4747_o;
  /* timer.vhd:227:9  */
  assign n4751_o = start_t_i ? 2'b01 : n4749_o;
  /* timer.vhd:194:7  */
  assign n4755_o = en_clk_i & n4737_o;
  /* timer.vhd:248:17  */
  assign n4773_o = read_timer_i ? counter_q : 8'b11111111;
  /* t48_pack-p.vhd:66:5  */
  assign n4782_o = overflow_q ? 1'b1 : 1'b0;
  /* timer.vhd:193:5  */
  assign n4783_o = en_clk_i ? n4728_o : counter_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4716_o)
    if (n4716_o)
      n4784_q <= 8'b00000000;
    else
      n4784_q <= n4783_o;
  /* timer.vhd:193:5  */
  assign n4785_o = en_clk_i ? n4730_o : overflow_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4716_o)
    if (n4716_o)
      n4786_q <= 1'b0;
    else
      n4786_q <= n4785_o;
  /* timer.vhd:193:5  */
  assign n4787_o = en_clk_i ? n4751_o : inc_sel_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4716_o)
    if (n4716_o)
      n4788_q <= 2'b00;
    else
      n4788_q <= n4787_o;
  /* timer.vhd:193:5  */
  assign n4789_o = n4755_o ? t1_i : t1_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4716_o)
    if (n4716_o)
      n4790_q <= 1'b0;
    else
      n4790_q <= n4789_o;
  /* timer.vhd:193:5  */
  assign n4791_o = en_clk_i ? n4745_o : prescaler_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4716_o)
    if (n4716_o)
      n4792_q <= 5'b00000;
    else
      n4792_q <= n4791_o;
endmodule

module t48_dmem_ctrl
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_dmem_addr_i,
   input  write_dmem_i,
   input  read_dmem_i,
   input  [1:0] addr_type_i,
   input  bank_select_i,
   input  [7:0] dmem_data_i,
   output [7:0] data_o,
   output [7:0] dmem_addr_o,
   output dmem_we_o,
   output [7:0] dmem_data_o);
  wire [7:0] dmem_addr_s;
  wire [7:0] dmem_addr_q;
  wire n4600_o;
  wire [2:0] n4601_o;
  localparam [7:0] n4602_o = 8'b00000000;
  wire [1:0] n4605_o;
  wire [1:0] n4606_o;
  wire [2:0] n4607_o;
  wire n4609_o;
  wire [2:0] n4610_o;
  wire [5:0] n4613_o;
  wire [5:0] n4615_o;
  localparam [7:0] n4616_o = 8'b00000000;
  wire [1:0] n4617_o;
  wire n4619_o;
  wire n4622_o;
  wire [3:0] n4623_o;
  wire n4624_o;
  wire n4625_o;
  wire n4626_o;
  wire n4627_o;
  reg n4628_o;
  wire [1:0] n4629_o;
  wire [1:0] n4630_o;
  wire [1:0] n4631_o;
  wire [1:0] n4632_o;
  reg [1:0] n4633_o;
  wire [1:0] n4634_o;
  wire [1:0] n4635_o;
  wire [1:0] n4636_o;
  reg [1:0] n4637_o;
  wire n4638_o;
  wire n4639_o;
  wire n4640_o;
  wire n4641_o;
  reg n4642_o;
  wire [1:0] n4643_o;
  wire [1:0] n4644_o;
  wire [1:0] n4645_o;
  reg [1:0] n4646_o;
  wire n4656_o;
  wire n4659_o;
  wire n4664_o;
  wire [7:0] n4665_o;
  wire [7:0] n4666_o;
  wire n4675_o;
  wire [7:0] n4676_o;
  wire [7:0] n4677_o;
  reg [7:0] n4678_q;
  assign data_o = n4666_o;
  assign dmem_addr_o = n4665_o;
  assign dmem_we_o = n4675_o;
  assign dmem_data_o = data_i;
  /* dmem_ctrl.vhd:91:10  */
  assign dmem_addr_s = n4676_o; // (signal)
  /* dmem_ctrl.vhd:92:10  */
  assign dmem_addr_q = n4678_q; // (signal)
  /* dmem_ctrl.vhd:112:7  */
  assign n4600_o = addr_type_i == 2'b00;
  /* dmem_ctrl.vhd:117:44  */
  assign n4601_o = data_i[2:0];
  /* decoder.vhd:155:5  */
  assign n4605_o = n4602_o[4:3];
  /* dmem_ctrl.vhd:119:9  */
  assign n4606_o = bank_select_i ? 2'b11 : n4605_o;
  /* decoder.vhd:153:5  */
  assign n4607_o = n4602_o[7:5];
  /* dmem_ctrl.vhd:115:7  */
  assign n4609_o = addr_type_i == 2'b01;
  /* dmem_ctrl.vhd:126:53  */
  assign n4610_o = data_i[2:0];
  /* decoder.vhd:142:5  */
  assign n4613_o = {2'b00, n4610_o, 1'b0};
  /* dmem_ctrl.vhd:128:51  */
  assign n4615_o = n4613_o + 6'b001000;
  /* decoder.vhd:135:5  */
  assign n4617_o = n4616_o[7:6];
  /* dmem_ctrl.vhd:124:7  */
  assign n4619_o = addr_type_i == 2'b10;
  /* dmem_ctrl.vhd:133:7  */
  assign n4622_o = addr_type_i == 2'b11;
  /* decoder.vhd:125:5  */
  assign n4623_o = {n4622_o, n4619_o, n4609_o, n4600_o};
  /* decoder.vhd:124:5  */
  assign n4624_o = data_i[0];
  /* decoder.vhd:123:5  */
  assign n4625_o = n4601_o[0];
  /* decoder.vhd:121:5  */
  assign n4626_o = n4615_o[0];
  /* decoder.vhd:120:5  */
  assign n4627_o = dmem_addr_q[0];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4623_o)
      4'b1000: n4628_o = 1'b1;
      4'b0100: n4628_o = n4626_o;
      4'b0010: n4628_o = n4625_o;
      4'b0001: n4628_o = n4624_o;
      default: n4628_o = n4627_o;
    endcase
  /* decoder.vhd:116:5  */
  assign n4629_o = data_i[2:1];
  /* decoder.vhd:115:5  */
  assign n4630_o = n4601_o[2:1];
  /* decoder.vhd:114:5  */
  assign n4631_o = n4615_o[2:1];
  /* decoder.vhd:113:5  */
  assign n4632_o = dmem_addr_q[2:1];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4623_o)
      4'b1000: n4633_o = n4632_o;
      4'b0100: n4633_o = n4631_o;
      4'b0010: n4633_o = n4630_o;
      4'b0001: n4633_o = n4629_o;
      default: n4633_o = n4632_o;
    endcase
  /* decoder.vhd:109:5  */
  assign n4634_o = data_i[4:3];
  /* decoder.vhd:108:5  */
  assign n4635_o = n4615_o[4:3];
  /* decoder.vhd:107:5  */
  assign n4636_o = dmem_addr_q[4:3];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4623_o)
      4'b1000: n4637_o = n4636_o;
      4'b0100: n4637_o = n4635_o;
      4'b0010: n4637_o = n4606_o;
      4'b0001: n4637_o = n4634_o;
      default: n4637_o = n4636_o;
    endcase
  /* decoder.vhd:105:5  */
  assign n4638_o = data_i[5];
  /* decoder.vhd:104:5  */
  assign n4639_o = n4607_o[0];
  /* decoder.vhd:103:5  */
  assign n4640_o = n4615_o[5];
  /* decoder.vhd:102:5  */
  assign n4641_o = dmem_addr_q[5];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4623_o)
      4'b1000: n4642_o = n4641_o;
      4'b0100: n4642_o = n4640_o;
      4'b0010: n4642_o = n4639_o;
      4'b0001: n4642_o = n4638_o;
      default: n4642_o = n4641_o;
    endcase
  /* decoder.vhd:100:5  */
  assign n4643_o = data_i[7:6];
  /* decoder.vhd:99:5  */
  assign n4644_o = n4607_o[2:1];
  /* decoder.vhd:98:5  */
  assign n4645_o = dmem_addr_q[7:6];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4623_o)
      4'b1000: n4646_o = n4645_o;
      4'b0100: n4646_o = n4617_o;
      4'b0010: n4646_o = n4644_o;
      4'b0001: n4646_o = n4643_o;
      default: n4646_o = n4645_o;
    endcase
  /* dmem_ctrl.vhd:165:14  */
  assign n4656_o = ~res_i;
  /* dmem_ctrl.vhd:169:7  */
  assign n4659_o = en_clk_i & write_dmem_addr_i;
  /* dmem_ctrl.vhd:188:41  */
  assign n4664_o = write_dmem_addr_i & en_clk_i;
  /* dmem_ctrl.vhd:188:18  */
  assign n4665_o = n4664_o ? dmem_addr_s : dmem_addr_q;
  /* dmem_ctrl.vhd:196:18  */
  assign n4666_o = read_dmem_i ? dmem_data_i : 8'b11111111;
  /* t48_pack-p.vhd:66:5  */
  assign n4675_o = write_dmem_i ? 1'b1 : 1'b0;
  assign n4676_o = {n4646_o, n4642_o, n4637_o, n4633_o, n4628_o};
  /* dmem_ctrl.vhd:168:5  */
  assign n4677_o = n4659_o ? dmem_addr_s : dmem_addr_q;
  /* dmem_ctrl.vhd:168:5  */
  always @(posedge clk_i or posedge n4656_o)
    if (n4656_o)
      n4678_q <= 8'b00000000;
    else
      n4678_q <= n4677_o;
endmodule

module t48_decoder_1_1_1
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  ea_i,
   input  ale_i,
   input  int_n_i,
   input  [7:0] data_i,
   input  bus_set_f1_i,
   input  bus_clear_f1_i,
   input  alu_carry_i,
   input  alu_da_overflow_i,
   input  [2:0] clk_mstate_i,
   input  clk_second_cycle_i,
   input  cnd_take_branch_i,
   input  psw_carry_i,
   input  psw_aux_carry_i,
   input  psw_f0_i,
   input  tim_overflow_i,
   output t0_dir_o,
   output [7:0] data_o,
   output alu_write_accu_o,
   output alu_write_shadow_o,
   output alu_write_temp_reg_o,
   output alu_read_alu_o,
   output bus_write_bus_o,
   output bus_read_bus_o,
   output bus_ibf_int_o,
   output bus_en_dma_o,
   output bus_en_flags_o,
   output bus_write_sts_o,
   output dm_write_dmem_addr_o,
   output dm_write_dmem_o,
   output dm_read_dmem_o,
   output p1_write_p1_o,
   output p1_read_p1_o,
   output p2_write_p2_o,
   output p2_write_exp_o,
   output p2_read_p2_o,
   output p2_read_exp_o,
   output pm_write_pcl_o,
   output pm_read_pcl_o,
   output pm_write_pch_o,
   output pm_read_pch_o,
   output pm_read_pmem_o,
   output psw_read_psw_o,
   output psw_read_sp_o,
   output psw_write_psw_o,
   output psw_write_sp_o,
   output [3:0] alu_op_o,
   output alu_use_carry_o,
   output alu_da_high_o,
   output alu_accu_low_o,
   output alu_p06_temp_reg_o,
   output alu_p60_temp_reg_o,
   output bus_output_pcl_o,
   output bus_bidir_bus_o,
   output clk_multi_cycle_o,
   output clk_assert_psen_o,
   output clk_assert_prog_o,
   output clk_assert_rd_o,
   output clk_assert_wr_o,
   output cnd_compute_take_o,
   output [3:0] cnd_branch_cond_o,
   output [2:0] cnd_comp_value_o,
   output cnd_f1_o,
   output cnd_tf_o,
   output [1:0] dm_addr_type_o,
   output p1_read_reg_o,
   output p2_read_reg_o,
   output p2_output_pch_o,
   output pm_inc_pc_o,
   output pm_write_pmem_addr_o,
   output [1:0] pm_addr_type_o,
   output psw_special_data_o,
   output psw_inc_stackp_o,
   output psw_dec_stackp_o,
   output psw_write_carry_o,
   output psw_write_aux_carry_o,
   output psw_write_f0_o,
   output psw_write_bs_o,
   output tim_read_timer_o,
   output tim_write_timer_o,
   output tim_start_t_o,
   output tim_start_cnt_o,
   output tim_stop_tcnt_o);
  wire opc_multi_cycle_s;
  wire opc_read_bus_s;
  wire opc_inj_int_s;
  wire [7:0] opc_opcode_q;
  wire [5:0] opc_mnemonic_s;
  wire last_cycle_s;
  wire assert_psen_s;
  wire branch_taken_s;
  wire branch_taken_q;
  wire pm_inc_pc_s;
  wire pm_write_pmem_addr_s;
  wire add_inc_pc_s;
  wire add_write_pmem_addr_s;
  wire clear_f1_s;
  wire cpl_f1_s;
  wire f1_q;
  wire clear_mb_s;
  wire set_mb_s;
  wire mb_q;
  wire ent0_clk_s;
  wire t0_dir_q;
  wire [7:0] data_s;
  wire read_dec_s;
  wire tf_s;
  wire bus_read_bus_s;
  wire add_read_bus_s;
  wire dm_write_dmem_s;
  wire p2_output_exp_s;
  wire movx_first_cycle_s;
  wire jtf_executed_s;
  wire en_tcnti_s;
  wire dis_tcnti_s;
  wire en_i_s;
  wire dis_i_s;
  wire tim_int_s;
  wire retr_executed_s;
  wire int_executed_s;
  wire int_pending_s;
  wire int_in_progress_s;
  wire [6:0] mnemonic_rec_s;
  wire [5:0] mnemonic_q;
  wire n1240_o;
  wire n1242_o;
  wire n1243_o;
  wire n1245_o;
  wire [1:0] n1246_o;
  reg [5:0] n1250_o;
  wire n1253_o;
  wire n1263_o;
  wire n1265_o;
  wire n1266_o;
  wire n1268_o;
  wire n1270_o;
  wire n1272_o;
  wire n1274_o;
  wire n1276_o;
  wire n1277_o;
  wire n1279_o;
  wire n1281_o;
  wire n1283_o;
  wire n1284_o;
  wire [6:0] n1285_o;
  reg [5:0] n1294_o;
  reg n1302_o;
  wire n1305_o;
  wire n1315_o;
  wire n1317_o;
  wire n1318_o;
  wire n1320_o;
  wire n1321_o;
  wire n1323_o;
  wire n1324_o;
  wire n1326_o;
  wire n1327_o;
  wire n1329_o;
  wire n1330_o;
  wire n1332_o;
  wire n1333_o;
  wire n1335_o;
  wire n1336_o;
  wire n1338_o;
  wire n1339_o;
  wire n1341_o;
  wire n1342_o;
  wire n1344_o;
  wire n1345_o;
  wire n1347_o;
  wire n1348_o;
  wire n1350_o;
  wire n1351_o;
  wire n1353_o;
  wire n1354_o;
  wire n1356_o;
  wire n1357_o;
  wire n1359_o;
  wire n1360_o;
  wire n1362_o;
  wire n1363_o;
  wire n1365_o;
  wire n1366_o;
  wire n1368_o;
  wire n1369_o;
  wire n1371_o;
  wire n1372_o;
  wire n1374_o;
  wire n1376_o;
  wire n1377_o;
  wire n1379_o;
  wire n1381_o;
  wire n1382_o;
  wire n1384_o;
  wire n1385_o;
  wire n1387_o;
  wire n1388_o;
  wire n1390_o;
  wire n1391_o;
  wire n1393_o;
  wire n1394_o;
  wire n1396_o;
  wire n1397_o;
  wire n1399_o;
  wire n1400_o;
  wire n1402_o;
  wire n1403_o;
  wire n1405_o;
  wire n1406_o;
  wire n1408_o;
  wire n1410_o;
  wire n1412_o;
  wire n1413_o;
  wire n1415_o;
  wire n1416_o;
  wire n1418_o;
  wire n1419_o;
  wire n1421_o;
  wire n1422_o;
  wire n1424_o;
  wire n1425_o;
  wire n1427_o;
  wire n1428_o;
  wire n1430_o;
  wire n1431_o;
  wire n1433_o;
  wire n1435_o;
  wire n1437_o;
  wire n1439_o;
  wire n1440_o;
  wire n1442_o;
  wire n1444_o;
  wire n1446_o;
  wire n1448_o;
  wire n1449_o;
  wire n1451_o;
  wire n1453_o;
  wire n1455_o;
  wire n1456_o;
  wire n1458_o;
  wire n1459_o;
  wire n1461_o;
  wire n1462_o;
  wire n1464_o;
  wire n1465_o;
  wire n1467_o;
  wire n1468_o;
  wire n1470_o;
  wire n1471_o;
  wire n1473_o;
  wire n1474_o;
  wire n1476_o;
  wire n1477_o;
  wire n1479_o;
  wire n1481_o;
  wire n1482_o;
  wire n1484_o;
  wire n1486_o;
  wire n1487_o;
  wire n1489_o;
  wire n1491_o;
  wire n1492_o;
  wire n1494_o;
  wire n1495_o;
  wire n1497_o;
  wire n1498_o;
  wire n1500_o;
  wire n1501_o;
  wire n1503_o;
  wire n1504_o;
  wire n1506_o;
  wire n1507_o;
  wire n1509_o;
  wire n1510_o;
  wire n1512_o;
  wire n1514_o;
  wire n1515_o;
  wire n1517_o;
  wire n1519_o;
  wire n1520_o;
  wire n1522_o;
  wire n1523_o;
  wire n1525_o;
  wire n1526_o;
  wire n1528_o;
  wire n1529_o;
  wire n1531_o;
  wire n1532_o;
  wire n1534_o;
  wire n1535_o;
  wire n1537_o;
  wire n1538_o;
  wire n1540_o;
  wire n1541_o;
  wire n1543_o;
  wire n1544_o;
  wire n1546_o;
  wire n1547_o;
  wire n1549_o;
  wire n1551_o;
  wire n1552_o;
  wire n1554_o;
  wire n1555_o;
  wire n1557_o;
  wire n1558_o;
  wire n1560_o;
  wire n1561_o;
  wire n1563_o;
  wire n1564_o;
  wire n1566_o;
  wire n1567_o;
  wire n1569_o;
  wire n1570_o;
  wire n1572_o;
  wire n1574_o;
  wire n1575_o;
  wire n1577_o;
  wire n1579_o;
  wire n1580_o;
  wire n1582_o;
  wire n1584_o;
  wire n1585_o;
  wire n1587_o;
  wire n1588_o;
  wire n1590_o;
  wire n1591_o;
  wire n1593_o;
  wire n1594_o;
  wire n1596_o;
  wire n1597_o;
  wire n1599_o;
  wire n1600_o;
  wire n1602_o;
  wire n1603_o;
  wire n1605_o;
  wire n1607_o;
  wire n1609_o;
  wire n1610_o;
  wire n1612_o;
  wire n1613_o;
  wire n1615_o;
  wire n1616_o;
  wire n1618_o;
  wire n1620_o;
  wire n1622_o;
  wire n1623_o;
  wire n1625_o;
  wire n1627_o;
  wire n1629_o;
  wire n1631_o;
  wire n1632_o;
  wire n1634_o;
  wire n1635_o;
  wire n1637_o;
  wire n1638_o;
  wire n1640_o;
  wire n1641_o;
  wire n1643_o;
  wire n1644_o;
  wire n1646_o;
  wire n1647_o;
  wire n1649_o;
  wire n1650_o;
  wire n1652_o;
  wire n1653_o;
  wire n1655_o;
  wire n1656_o;
  wire n1658_o;
  wire n1660_o;
  wire n1662_o;
  wire n1663_o;
  wire n1665_o;
  wire n1666_o;
  wire n1668_o;
  wire n1669_o;
  wire n1671_o;
  wire n1672_o;
  wire n1674_o;
  wire n1675_o;
  wire n1677_o;
  wire n1678_o;
  wire n1680_o;
  wire n1681_o;
  wire n1683_o;
  wire n1684_o;
  wire n1686_o;
  wire n1687_o;
  wire n1689_o;
  wire n1691_o;
  wire n1692_o;
  wire n1694_o;
  wire n1695_o;
  wire n1697_o;
  wire n1698_o;
  wire n1700_o;
  wire n1701_o;
  wire n1703_o;
  wire n1704_o;
  wire n1706_o;
  wire n1707_o;
  wire n1709_o;
  wire n1710_o;
  wire n1712_o;
  wire n1713_o;
  wire n1715_o;
  wire n1716_o;
  wire n1718_o;
  wire n1720_o;
  wire n1721_o;
  wire n1723_o;
  wire n1725_o;
  wire n1726_o;
  wire n1728_o;
  wire n1729_o;
  wire n1731_o;
  wire n1732_o;
  wire n1734_o;
  wire n1736_o;
  wire n1737_o;
  wire n1739_o;
  wire n1741_o;
  wire n1743_o;
  wire n1744_o;
  wire n1746_o;
  wire n1747_o;
  wire n1749_o;
  wire n1750_o;
  wire n1752_o;
  wire n1753_o;
  wire n1755_o;
  wire n1756_o;
  wire n1758_o;
  wire n1759_o;
  wire n1761_o;
  wire n1762_o;
  wire n1764_o;
  wire n1765_o;
  wire n1767_o;
  wire n1768_o;
  wire n1770_o;
  wire n1772_o;
  wire n1774_o;
  wire n1775_o;
  wire n1777_o;
  wire n1778_o;
  wire n1780_o;
  wire n1781_o;
  wire n1783_o;
  wire n1784_o;
  wire n1786_o;
  wire n1787_o;
  wire n1789_o;
  wire n1790_o;
  wire n1792_o;
  wire n1793_o;
  wire n1795_o;
  wire n1796_o;
  wire n1798_o;
  wire n1799_o;
  wire n1801_o;
  wire n1802_o;
  wire n1804_o;
  wire n1805_o;
  wire n1807_o;
  wire n1809_o;
  wire n1810_o;
  wire n1812_o;
  wire n1814_o;
  wire n1815_o;
  wire n1817_o;
  wire n1819_o;
  wire n1820_o;
  wire n1822_o;
  wire n1824_o;
  wire n1825_o;
  wire n1827_o;
  wire n1829_o;
  wire n1831_o;
  wire n1832_o;
  wire n1834_o;
  wire n1836_o;
  wire n1838_o;
  wire n1839_o;
  wire n1841_o;
  wire n1842_o;
  wire n1844_o;
  wire n1845_o;
  wire n1847_o;
  wire n1848_o;
  wire n1850_o;
  wire n1851_o;
  wire n1853_o;
  wire n1854_o;
  wire n1856_o;
  wire n1857_o;
  wire n1859_o;
  wire n1860_o;
  wire n1862_o;
  wire n1863_o;
  wire n1865_o;
  wire n1866_o;
  wire n1868_o;
  wire n1869_o;
  wire n1871_o;
  wire n1873_o;
  wire n1874_o;
  wire n1876_o;
  wire n1877_o;
  wire n1879_o;
  wire n1880_o;
  wire n1882_o;
  wire n1883_o;
  wire n1885_o;
  wire n1886_o;
  wire n1888_o;
  wire n1889_o;
  wire n1891_o;
  wire n1892_o;
  wire n1894_o;
  wire n1895_o;
  wire n1897_o;
  wire n1898_o;
  wire n1900_o;
  wire [48:0] n1901_o;
  reg [5:0] n1952_o;
  reg n1976_o;
  wire [6:0] n1980_o;
  wire [6:0] n1981_o;
  wire [6:0] n1982_o;
  wire [6:0] n1985_o;
  wire [6:0] n1986_o;
  wire n1989_o;
  wire [5:0] n1991_o;
  wire [7:0] n1993_o;
  wire [5:0] n1994_o;
  wire [7:0] n1995_o;
  wire [5:0] n1996_o;
  wire n2006_o;
  wire [5:0] n2008_o;
  wire [5:0] n2009_o;
  wire int_b_n2010;
  wire int_b_n2012;
  wire int_b_n2013;
  wire int_b_n2014;
  wire int_b_tf_o;
  wire int_b_ext_int_o;
  wire int_b_tim_int_o;
  wire int_b_int_pending_o;
  wire int_b_int_in_progress_o;
  wire n2024_o;
  wire n2025_o;
  wire n2026_o;
  wire n2029_o;
  wire n2030_o;
  wire n2031_o;
  wire n2032_o;
  wire n2033_o;
  wire n2036_o;
  wire n2037_o;
  wire n2040_o;
  wire n2042_o;
  wire n2045_o;
  wire n2047_o;
  wire n2049_o;
  wire n2051_o;
  wire n2053_o;
  wire n2054_o;
  wire n2055_o;
  wire n2058_o;
  wire n2061_o;
  wire n2063_o;
  wire n2065_o;
  wire n2067_o;
  wire n2068_o;
  wire n2069_o;
  wire n2070_o;
  wire n2071_o;
  wire n2074_o;
  wire n2076_o;
  wire n2079_o;
  wire n2081_o;
  wire n2082_o;
  wire n2083_o;
  wire n2084_o;
  wire n2085_o;
  wire n2088_o;
  wire n2091_o;
  wire n2094_o;
  wire n2096_o;
  wire n2097_o;
  wire n2098_o;
  wire n2099_o;
  wire n2100_o;
  wire n2101_o;
  wire n2102_o;
  wire n2105_o;
  wire n2107_o;
  wire [4:0] n2108_o;
  reg n2110_o;
  reg n2113_o;
  reg n2116_o;
  reg n2119_o;
  reg n2122_o;
  reg n2125_o;
  reg n2128_o;
  reg n2131_o;
  reg n2134_o;
  wire n2141_o;
  wire n2142_o;
  wire n2144_o;
  wire n2145_o;
  wire n2146_o;
  wire [2:0] n2147_o;
  wire n2148_o;
  wire [2:0] n2150_o;
  wire [2:0] n2151_o;
  localparam [7:0] n2152_o = 8'b00000000;
  wire [4:0] n2153_o;
  wire n2156_o;
  wire [7:0] n2158_o;
  localparam [7:0] n2159_o = 8'bX;
  wire [7:0] n2160_o;
  wire n2164_o;
  wire n2166_o;
  wire n2167_o;
  wire n2169_o;
  wire n2176_o;
  wire n2179_o;
  wire [1:0] n2182_o;
  wire n2184_o;
  wire n2189_o;
  wire n2193_o;
  wire n2196_o;
  wire n2198_o;
  wire [2:0] n2199_o;
  reg n2202_o;
  reg n2205_o;
  reg n2208_o;
  reg n2209_o;
  reg n2212_o;
  reg [3:0] n2215_o;
  reg n2217_o;
  reg [1:0] n2219_o;
  reg n2221_o;
  reg n2224_o;
  reg n2227_o;
  wire n2229_o;
  wire n2231_o;
  wire n2235_o;
  wire n2238_o;
  wire n2240_o;
  wire [1:0] n2241_o;
  reg n2244_o;
  reg n2247_o;
  reg n2250_o;
  reg [3:0] n2253_o;
  reg n2255_o;
  reg n2257_o;
  reg n2260_o;
  reg n2263_o;
  wire n2265_o;
  wire n2267_o;
  wire n2269_o;
  wire [3:0] n2271_o;
  wire n2273_o;
  wire n2275_o;
  wire n2277_o;
  wire n2279_o;
  wire n2281_o;
  wire n2282_o;
  wire n2283_o;
  wire n2285_o;
  wire n2292_o;
  wire n2295_o;
  wire [1:0] n2298_o;
  wire n2300_o;
  wire n2305_o;
  wire n2310_o;
  wire [2:0] n2311_o;
  reg n2314_o;
  reg n2317_o;
  reg n2320_o;
  reg n2321_o;
  reg n2324_o;
  reg [3:0] n2327_o;
  reg [1:0] n2329_o;
  wire n2331_o;
  wire n2333_o;
  wire n2338_o;
  wire [1:0] n2339_o;
  reg n2342_o;
  reg n2345_o;
  reg n2348_o;
  reg [3:0] n2351_o;
  wire n2353_o;
  wire n2355_o;
  wire n2357_o;
  wire [3:0] n2359_o;
  wire n2361_o;
  wire n2362_o;
  wire n2364_o;
  wire [1:0] n2365_o;
  wire n2367_o;
  wire n2368_o;
  wire n2369_o;
  wire n2372_o;
  wire n2375_o;
  wire n2378_o;
  wire n2381_o;
  wire n2383_o;
  wire n2385_o;
  wire n2387_o;
  wire n2389_o;
  wire n2392_o;
  wire n2395_o;
  wire n2397_o;
  wire n2399_o;
  wire n2401_o;
  wire n2403_o;
  wire n2405_o;
  wire n2407_o;
  wire n2409_o;
  wire [1:0] n2410_o;
  wire n2412_o;
  wire n2413_o;
  wire n2414_o;
  wire n2417_o;
  wire n2420_o;
  wire n2423_o;
  wire n2425_o;
  wire n2427_o;
  wire n2429_o;
  wire [2:0] n2430_o;
  reg n2434_o;
  reg n2438_o;
  reg n2440_o;
  reg n2442_o;
  reg n2444_o;
  reg [3:0] n2447_o;
  wire n2449_o;
  wire n2451_o;
  wire n2453_o;
  wire n2455_o;
  wire n2457_o;
  wire n2459_o;
  wire n2461_o;
  wire n2463_o;
  wire [3:0] n2465_o;
  wire n2467_o;
  wire n2469_o;
  wire n2471_o;
  wire n2473_o;
  wire n2474_o;
  wire n2475_o;
  wire n2478_o;
  wire n2480_o;
  wire n2482_o;
  wire n2484_o;
  wire [2:0] n2485_o;
  reg n2488_o;
  reg n2491_o;
  reg n2494_o;
  reg n2497_o;
  reg n2500_o;
  reg [1:0] n2504_o;
  reg n2507_o;
  reg n2509_o;
  reg n2513_o;
  localparam [7:0] n2515_o = 8'b00000000;
  wire n2520_o;
  wire n2521_o;
  wire n2522_o;
  wire [4:0] n2523_o;
  wire n2525_o;
  wire [7:0] n2526_o;
  wire [7:0] n2527_o;
  wire n2529_o;
  wire n2531_o;
  wire n2532_o;
  wire [4:0] n2534_o;
  wire [2:0] n2535_o;
  wire [7:0] n2536_o;
  wire [7:0] n2538_o;
  wire n2541_o;
  wire n2543_o;
  wire [1:0] n2544_o;
  reg n2546_o;
  reg n2549_o;
  reg n2552_o;
  reg n2555_o;
  reg [7:0] n2556_o;
  reg n2558_o;
  reg n2560_o;
  wire n2562_o;
  wire n2563_o;
  wire n2565_o;
  wire n2567_o;
  wire n2569_o;
  wire n2571_o;
  wire n2573_o;
  wire n2575_o;
  wire [1:0] n2577_o;
  wire n2579_o;
  wire n2581_o;
  wire n2583_o;
  wire [7:0] n2584_o;
  wire n2585_o;
  wire n2587_o;
  wire n2589_o;
  wire n2591_o;
  wire n2593_o;
  wire n2596_o;
  wire n2599_o;
  wire [3:0] n2602_o;
  wire n2604_o;
  wire n2606_o;
  wire n2609_o;
  wire n2611_o;
  wire n2613_o;
  wire n2614_o;
  wire n2615_o;
  wire n2618_o;
  wire n2621_o;
  wire n2623_o;
  wire n2625_o;
  wire n2627_o;
  wire n2629_o;
  wire n2632_o;
  wire n2635_o;
  wire [3:0] n2638_o;
  wire n2640_o;
  wire n2642_o;
  wire n2643_o;
  wire n2645_o;
  wire n2648_o;
  wire n2650_o;
  wire n2652_o;
  wire n2653_o;
  wire n2654_o;
  wire n2655_o;
  wire n2657_o;
  wire n2660_o;
  wire n2663_o;
  wire n2665_o;
  wire n2667_o;
  wire n2669_o;
  wire n2671_o;
  wire n2673_o;
  wire n2674_o;
  wire n2677_o;
  wire n2680_o;
  wire n2682_o;
  wire [3:0] n2685_o;
  wire n2687_o;
  wire n2689_o;
  wire [2:0] n2690_o;
  reg n2693_o;
  reg n2695_o;
  reg n2698_o;
  reg [3:0] n2700_o;
  reg n2704_o;
  reg n2707_o;
  reg n2710_o;
  reg n2712_o;
  reg n2715_o;
  wire n2717_o;
  wire n2718_o;
  wire n2721_o;
  wire n2724_o;
  wire n2726_o;
  wire n2727_o;
  wire n2728_o;
  wire n2731_o;
  wire n2734_o;
  wire n2736_o;
  wire [1:0] n2737_o;
  reg n2739_o;
  reg n2741_o;
  reg n2744_o;
  reg n2746_o;
  reg [3:0] n2749_o;
  reg n2751_o;
  wire n2753_o;
  wire n2755_o;
  wire n2756_o;
  wire n2759_o;
  wire n2762_o;
  wire n2764_o;
  wire n2766_o;
  wire n2768_o;
  wire n2770_o;
  wire n2771_o;
  wire n2774_o;
  wire n2777_o;
  wire n2779_o;
  wire n2781_o;
  wire n2783_o;
  wire n2784_o;
  wire n2786_o;
  wire n2789_o;
  wire [1:0] n2790_o;
  reg n2793_o;
  reg n2796_o;
  reg n2799_o;
  reg [3:0] n2802_o;
  reg n2805_o;
  reg [3:0] n2808_o;
  wire n2809_o;
  reg n2810_o;
  reg n2813_o;
  wire n2815_o;
  wire n2816_o;
  wire n2822_o;
  wire n2825_o;
  wire n2827_o;
  wire n2829_o;
  wire n2831_o;
  wire n2833_o;
  wire [3:0] n2835_o;
  wire n2837_o;
  wire [3:0] n2839_o;
  wire n2840_o;
  wire n2841_o;
  wire n2843_o;
  wire n2845_o;
  wire n2847_o;
  wire n2849_o;
  wire n2850_o;
  wire n2851_o;
  wire n2854_o;
  wire n2857_o;
  wire n2859_o;
  wire n2861_o;
  wire n2863_o;
  wire n2865_o;
  wire n2868_o;
  wire n2870_o;
  wire n2872_o;
  wire n2873_o;
  wire n2874_o;
  wire n2875_o;
  wire n2878_o;
  wire n2881_o;
  wire n2884_o;
  wire n2886_o;
  wire n2888_o;
  wire n2890_o;
  wire n2892_o;
  wire n2895_o;
  wire n2898_o;
  wire n2900_o;
  wire n2902_o;
  wire n2903_o;
  wire n2906_o;
  wire n2909_o;
  wire n2911_o;
  wire n2912_o;
  wire n2913_o;
  wire n2915_o;
  wire n2922_o;
  wire n2925_o;
  wire [1:0] n2928_o;
  wire n2930_o;
  wire [1:0] n2931_o;
  wire n2933_o;
  wire n2936_o;
  wire n2939_o;
  wire n2941_o;
  wire [1:0] n2942_o;
  wire n2944_o;
  wire n2947_o;
  wire n2950_o;
  wire n2952_o;
  wire [2:0] n2953_o;
  reg n2955_o;
  reg n2957_o;
  reg n2960_o;
  reg n2961_o;
  reg n2963_o;
  reg [3:0] n2966_o;
  reg [1:0] n2968_o;
  reg n2970_o;
  wire n2972_o;
  wire n2973_o;
  wire n2975_o;
  wire n2978_o;
  wire n2981_o;
  wire n2983_o;
  wire n2984_o;
  wire n2990_o;
  wire n2993_o;
  wire n2995_o;
  wire n2997_o;
  wire n2999_o;
  wire n3001_o;
  wire n3003_o;
  wire n3004_o;
  wire n3006_o;
  wire n3007_o;
  wire n3010_o;
  wire n3011_o;
  wire n3012_o;
  wire n3014_o;
  wire n3015_o;
  wire n3021_o;
  wire n3024_o;
  wire n3026_o;
  wire n3028_o;
  wire n3030_o;
  wire n3032_o;
  wire n3034_o;
  wire n3035_o;
  wire n3037_o;
  wire n3038_o;
  wire [3:0] n3041_o;
  wire n3044_o;
  wire [3:0] n3046_o;
  wire n3048_o;
  wire n3049_o;
  wire n3055_o;
  wire n3058_o;
  wire n3060_o;
  wire n3062_o;
  wire [3:0] n3064_o;
  wire n3066_o;
  wire n3068_o;
  wire n3070_o;
  wire [4:0] n3072_o;
  wire [2:0] n3073_o;
  wire [7:0] n3074_o;
  wire n3076_o;
  wire [1:0] n3077_o;
  reg n3080_o;
  reg n3083_o;
  reg n3086_o;
  reg [7:0] n3087_o;
  reg n3089_o;
  wire n3091_o;
  wire n3093_o;
  wire n3095_o;
  wire [7:0] n3096_o;
  wire n3097_o;
  wire n3099_o;
  wire n3100_o;
  wire n3102_o;
  wire n3105_o;
  wire [1:0] n3108_o;
  wire n3110_o;
  wire n3113_o;
  wire n3116_o;
  wire n3118_o;
  wire n3120_o;
  wire [1:0] n3122_o;
  wire n3124_o;
  wire n3126_o;
  wire n3127_o;
  wire n3129_o;
  wire n3132_o;
  wire n3134_o;
  wire n3135_o;
  wire n3141_o;
  wire n3144_o;
  wire n3146_o;
  wire n3148_o;
  wire n3150_o;
  wire n3152_o;
  wire n3153_o;
  wire n3155_o;
  wire n3158_o;
  wire n3160_o;
  wire n3161_o;
  wire n3167_o;
  wire n3170_o;
  wire n3172_o;
  wire n3174_o;
  wire n3176_o;
  wire n3178_o;
  wire n3179_o;
  wire n3181_o;
  wire n3184_o;
  wire n3186_o;
  wire n3187_o;
  wire n3193_o;
  wire n3196_o;
  wire n3198_o;
  wire n3200_o;
  wire n3202_o;
  wire n3204_o;
  wire n3205_o;
  wire n3206_o;
  wire [3:0] n3209_o;
  wire n3210_o;
  wire n3212_o;
  wire n3213_o;
  wire n3216_o;
  wire n3217_o;
  wire n3218_o;
  wire n3220_o;
  wire n3221_o;
  wire n3227_o;
  wire n3230_o;
  wire n3232_o;
  wire n3234_o;
  wire n3236_o;
  wire n3238_o;
  wire n3240_o;
  wire n3241_o;
  wire n3243_o;
  wire n3246_o;
  wire n3249_o;
  wire n3251_o;
  wire n3252_o;
  wire n3258_o;
  wire n3261_o;
  wire n3263_o;
  wire n3265_o;
  wire n3267_o;
  wire n3269_o;
  wire n3271_o;
  wire n3272_o;
  wire n3274_o;
  wire n3275_o;
  wire n3278_o;
  wire n3281_o;
  wire n3282_o;
  wire n3283_o;
  wire n3285_o;
  wire n3286_o;
  wire n3292_o;
  wire n3295_o;
  wire n3297_o;
  wire n3299_o;
  wire n3301_o;
  wire n3303_o;
  wire n3305_o;
  wire n3307_o;
  wire n3309_o;
  wire n3310_o;
  wire n3313_o;
  wire n3315_o;
  wire n3316_o;
  wire n3317_o;
  wire n3319_o;
  wire n3326_o;
  wire n3329_o;
  wire [1:0] n3332_o;
  wire n3334_o;
  wire n3339_o;
  wire [1:0] n3340_o;
  reg n3343_o;
  reg n3346_o;
  reg n3347_o;
  reg n3350_o;
  reg [1:0] n3352_o;
  wire n3354_o;
  wire n3356_o;
  wire n3359_o;
  wire n3362_o;
  wire n3365_o;
  wire n3367_o;
  wire n3369_o;
  wire n3372_o;
  wire n3375_o;
  wire n3378_o;
  wire n3380_o;
  wire n3381_o;
  wire n3382_o;
  wire n3384_o;
  wire n3391_o;
  wire n3394_o;
  wire [1:0] n3397_o;
  wire n3399_o;
  wire n3401_o;
  wire [1:0] n3402_o;
  reg n3405_o;
  reg n3406_o;
  reg n3408_o;
  reg [1:0] n3410_o;
  reg n3413_o;
  wire n3415_o;
  wire n3416_o;
  wire n3418_o;
  wire n3419_o;
  wire n3420_o;
  wire n3421_o;
  wire n3423_o;
  wire n3430_o;
  wire n3433_o;
  wire [1:0] n3436_o;
  wire n3437_o;
  wire n3439_o;
  wire [1:0] n3441_o;
  wire n3443_o;
  wire n3444_o;
  wire n3447_o;
  wire n3449_o;
  wire n3451_o;
  wire n3454_o;
  wire n3457_o;
  wire n3459_o;
  wire n3461_o;
  wire n3462_o;
  wire n3465_o;
  wire n3468_o;
  wire n3471_o;
  wire n3474_o;
  wire n3476_o;
  wire n3478_o;
  wire n3480_o;
  wire n3482_o;
  wire n3484_o;
  wire n3485_o;
  wire [1:0] n3487_o;
  wire [3:0] n3488_o;
  wire n3491_o;
  wire n3494_o;
  wire n3497_o;
  wire [2:0] n3498_o;
  wire [1:0] n3499_o;
  wire [1:0] n3500_o;
  wire [1:0] n3501_o;
  reg [1:0] n3502_o;
  wire n3504_o;
  wire n3506_o;
  wire n3508_o;
  wire [2:0] n3509_o;
  reg n3512_o;
  reg n3516_o;
  wire [1:0] n3517_o;
  wire [1:0] n3518_o;
  wire [1:0] n3519_o;
  reg [1:0] n3520_o;
  wire [1:0] n3521_o;
  wire [1:0] n3522_o;
  wire [1:0] n3523_o;
  reg [1:0] n3524_o;
  wire [3:0] n3525_o;
  wire [3:0] n3526_o;
  wire [3:0] n3527_o;
  reg [3:0] n3528_o;
  reg n3530_o;
  reg n3534_o;
  wire n3536_o;
  wire n3538_o;
  wire n3539_o;
  wire n3542_o;
  wire n3544_o;
  wire n3546_o;
  wire [7:0] n3547_o;
  wire [7:0] n3548_o;
  wire n3549_o;
  wire n3550_o;
  wire n3552_o;
  wire n3553_o;
  wire [1:0] n3554_o;
  wire [7:0] n3556_o;
  wire n3558_o;
  wire n3561_o;
  wire n3563_o;
  wire [2:0] n3564_o;
  reg n3568_o;
  wire [3:0] n3569_o;
  wire [3:0] n3570_o;
  wire [3:0] n3571_o;
  wire [3:0] n3572_o;
  reg [3:0] n3573_o;
  wire [3:0] n3574_o;
  wire [3:0] n3575_o;
  wire [3:0] n3576_o;
  wire [3:0] n3577_o;
  reg [3:0] n3578_o;
  reg n3581_o;
  reg n3585_o;
  wire n3587_o;
  wire n3589_o;
  wire [1:0] n3590_o;
  reg n3593_o;
  reg n3596_o;
  reg n3599_o;
  reg n3603_o;
  wire n3605_o;
  wire n3607_o;
  wire n3609_o;
  wire n3611_o;
  wire [7:0] n3612_o;
  wire [7:0] n3613_o;
  wire n3614_o;
  wire n3615_o;
  wire n3617_o;
  wire n3618_o;
  wire n3620_o;
  wire n3621_o;
  wire n3622_o;
  wire [1:0] n3625_o;
  wire n3628_o;
  wire [1:0] n3630_o;
  wire n3632_o;
  wire n3635_o;
  wire n3638_o;
  wire n3640_o;
  wire n3642_o;
  wire [1:0] n3644_o;
  wire n3646_o;
  wire n3648_o;
  wire n3649_o;
  wire n3650_o;
  wire n3653_o;
  wire n3656_o;
  wire n3657_o;
  wire n3659_o;
  wire n3660_o;
  wire n3663_o;
  wire n3666_o;
  wire n3668_o;
  wire [1:0] n3669_o;
  reg n3671_o;
  reg n3674_o;
  reg n3677_o;
  wire n3679_o;
  wire n3680_o;
  wire n3681_o;
  wire n3684_o;
  wire n3687_o;
  wire n3690_o;
  wire n3693_o;
  wire n3695_o;
  wire n3697_o;
  wire n3699_o;
  wire n3701_o;
  wire n3703_o;
  wire n3704_o;
  wire n3705_o;
  wire n3707_o;
  wire n3709_o;
  wire n3712_o;
  wire n3714_o;
  wire n3716_o;
  wire n3717_o;
  wire n3718_o;
  wire n3720_o;
  wire n3727_o;
  wire n3730_o;
  wire [1:0] n3733_o;
  wire n3735_o;
  wire n3740_o;
  wire n3745_o;
  wire [2:0] n3746_o;
  reg n3749_o;
  reg n3752_o;
  reg n3755_o;
  reg n3756_o;
  reg n3759_o;
  reg [3:0] n3762_o;
  reg [1:0] n3764_o;
  wire n3766_o;
  wire n3768_o;
  wire n3773_o;
  wire [1:0] n3774_o;
  reg n3777_o;
  reg n3780_o;
  reg n3783_o;
  reg [3:0] n3786_o;
  wire n3788_o;
  wire n3790_o;
  wire n3792_o;
  wire [3:0] n3794_o;
  wire n3796_o;
  wire n3797_o;
  wire n3799_o;
  wire [1:0] n3800_o;
  wire n3802_o;
  wire n3803_o;
  wire n3804_o;
  wire n3807_o;
  wire n3810_o;
  wire n3813_o;
  wire n3816_o;
  wire n3818_o;
  wire n3820_o;
  wire n3822_o;
  wire n3824_o;
  wire n3827_o;
  wire n3830_o;
  wire n3832_o;
  wire n3834_o;
  wire n3836_o;
  wire n3838_o;
  wire n3840_o;
  wire n3842_o;
  wire n3844_o;
  wire [1:0] n3845_o;
  wire n3847_o;
  wire n3848_o;
  wire n3849_o;
  wire n3852_o;
  wire n3855_o;
  wire n3858_o;
  wire n3860_o;
  wire n3862_o;
  wire n3864_o;
  wire [2:0] n3865_o;
  reg n3869_o;
  reg n3873_o;
  reg n3875_o;
  reg n3877_o;
  reg n3879_o;
  reg [3:0] n3882_o;
  wire n3884_o;
  wire n3886_o;
  wire n3888_o;
  wire n3890_o;
  wire n3892_o;
  wire n3894_o;
  wire n3896_o;
  wire n3898_o;
  wire [3:0] n3900_o;
  wire n3902_o;
  wire n3904_o;
  wire n3906_o;
  wire n3908_o;
  wire n3910_o;
  wire n3913_o;
  wire n3916_o;
  wire n3918_o;
  wire n3919_o;
  wire n3920_o;
  wire n3923_o;
  wire n3924_o;
  wire n3926_o;
  wire n3927_o;
  wire n3928_o;
  wire n3929_o;
  wire n3930_o;
  wire n3933_o;
  wire n3936_o;
  wire n3939_o;
  wire n3941_o;
  wire n3943_o;
  wire n3946_o;
  wire n3948_o;
  wire n3950_o;
  wire n3952_o;
  wire n3954_o;
  wire n3955_o;
  wire n3957_o;
  wire n3959_o;
  wire n3961_o;
  wire [2:0] n3962_o;
  reg n3965_o;
  reg n3968_o;
  reg n3971_o;
  reg n3974_o;
  reg [1:0] n3978_o;
  reg n3981_o;
  wire n3982_o;
  wire n3985_o;
  wire n3988_o;
  wire n3990_o;
  wire n3992_o;
  wire [1:0] n3993_o;
  reg n3996_o;
  reg n3999_o;
  reg n4001_o;
  reg n4004_o;
  reg n4006_o;
  wire n4007_o;
  wire n4008_o;
  wire n4010_o;
  wire n4012_o;
  wire n4014_o;
  wire n4016_o;
  wire [1:0] n4018_o;
  wire n4020_o;
  wire n4022_o;
  wire n4024_o;
  wire n4026_o;
  wire n4028_o;
  wire n4029_o;
  wire n4032_o;
  wire n4034_o;
  wire n4037_o;
  wire n4040_o;
  wire n4043_o;
  wire [3:0] n4046_o;
  wire n4048_o;
  wire n4050_o;
  wire n4052_o;
  wire n4054_o;
  wire n4056_o;
  wire n4057_o;
  wire n4058_o;
  wire n4061_o;
  wire n4063_o;
  wire n4066_o;
  wire n4069_o;
  wire n4072_o;
  wire [3:0] n4075_o;
  wire n4077_o;
  wire n4079_o;
  wire n4081_o;
  wire n4083_o;
  wire n4085_o;
  wire n4086_o;
  wire n4089_o;
  wire n4092_o;
  wire n4094_o;
  wire n4096_o;
  wire n4098_o;
  wire n4100_o;
  wire n4101_o;
  wire n4103_o;
  wire n4106_o;
  wire n4108_o;
  wire n4110_o;
  wire n4113_o;
  wire n4115_o;
  wire n4117_o;
  wire n4118_o;
  wire n4121_o;
  wire n4124_o;
  wire n4126_o;
  wire n4128_o;
  wire n4130_o;
  wire n4132_o;
  wire n4135_o;
  wire n4138_o;
  wire n4140_o;
  wire n4141_o;
  wire n4142_o;
  wire n4144_o;
  wire n4151_o;
  wire n4154_o;
  wire [1:0] n4157_o;
  wire n4159_o;
  wire n4160_o;
  wire n4163_o;
  wire n4165_o;
  wire n4166_o;
  wire [3:0] n4169_o;
  wire n4171_o;
  wire [2:0] n4172_o;
  reg n4175_o;
  reg n4178_o;
  reg n4181_o;
  reg n4182_o;
  reg n4185_o;
  reg [3:0] n4187_o;
  reg n4189_o;
  reg [1:0] n4191_o;
  reg n4194_o;
  wire n4196_o;
  wire n4197_o;
  wire n4198_o;
  wire n4200_o;
  wire n4207_o;
  wire n4210_o;
  wire [1:0] n4213_o;
  wire n4215_o;
  wire n4220_o;
  wire n4225_o;
  wire [2:0] n4226_o;
  reg n4229_o;
  reg n4232_o;
  reg n4235_o;
  reg n4236_o;
  reg n4239_o;
  reg [3:0] n4242_o;
  reg [1:0] n4244_o;
  wire n4246_o;
  wire n4248_o;
  wire n4253_o;
  wire [1:0] n4254_o;
  reg n4257_o;
  reg n4260_o;
  reg n4263_o;
  reg [3:0] n4266_o;
  wire n4268_o;
  wire n4270_o;
  wire n4272_o;
  wire [3:0] n4274_o;
  wire n4276_o;
  wire [62:0] n4277_o;
  reg n4279_o;
  reg n4282_o;
  reg n4285_o;
  reg n4288_o;
  reg n4291_o;
  reg n4294_o;
  reg n4297_o;
  reg n4300_o;
  reg n4303_o;
  reg n4305_o;
  reg n4307_o;
  reg n4310_o;
  reg n4313_o;
  reg n4316_o;
  reg n4319_o;
  reg n4322_o;
  reg n4325_o;
  reg n4328_o;
  reg n4331_o;
  reg n4334_o;
  reg n4337_o;
  reg n4340_o;
  reg n4343_o;
  reg n4346_o;
  reg n4349_o;
  reg [3:0] n4353_o;
  reg n4356_o;
  reg n4359_o;
  reg n4362_o;
  reg n4365_o;
  reg n4368_o;
  reg n4372_o;
  reg n4377_o;
  reg n4381_o;
  reg n4384_o;
  reg n4387_o;
  reg [3:0] n4397_o;
  wire n4399_o;
  reg n4400_o;
  wire [1:0] n4401_o;
  reg [1:0] n4403_o;
  reg n4406_o;
  reg n4409_o;
  reg [1:0] n4412_o;
  reg n4415_o;
  reg n4418_o;
  reg n4421_o;
  reg n4424_o;
  reg n4427_o;
  reg n4430_o;
  reg n4433_o;
  reg n4436_o;
  reg n4439_o;
  reg n4442_o;
  reg n4445_o;
  reg n4448_o;
  reg n4473_o;
  reg n4476_o;
  reg n4479_o;
  reg n4482_o;
  reg n4485_o;
  reg n4488_o;
  reg n4491_o;
  reg n4494_o;
  reg n4497_o;
  reg [7:0] n4499_o;
  reg n4500_o;
  reg n4502_o;
  reg n4505_o;
  reg n4508_o;
  reg n4511_o;
  reg n4514_o;
  reg n4517_o;
  reg n4520_o;
  reg n4523_o;
  reg n4526_o;
  reg n4529_o;
  reg n4532_o;
  wire n4536_o;
  wire n4539_o;
  wire n4541_o;
  wire n4543_o;
  wire n4545_o;
  wire n4547_o;
  wire n4548_o;
  wire n4549_o;
  wire n4551_o;
  wire n4553_o;
  wire n4555_o;
  wire n4559_o;
  wire n4561_o;
  wire [7:0] n4575_o;
  wire n4577_o;
  wire n4578_o;
  wire n4579_o;
  wire n4580_o;
  wire [7:0] n4581_o;
  reg [7:0] n4582_q;
  wire n4583_o;
  reg n4584_q;
  reg n4585_q;
  wire n4586_o;
  reg n4587_q;
  wire n4588_o;
  reg n4589_q;
  wire [5:0] n4590_o;
  reg [5:0] n4591_q;
  wire [2:0] n4592_o;
  assign t0_dir_o = t0_dir_q;
  assign data_o = n4575_o;
  assign alu_write_accu_o = n4279_o;
  assign alu_write_shadow_o = n4282_o;
  assign alu_write_temp_reg_o = n4285_o;
  assign alu_read_alu_o = n4288_o;
  assign bus_write_bus_o = n4291_o;
  assign bus_read_bus_o = n4580_o;
  assign bus_ibf_int_o = n4294_o;
  assign bus_en_dma_o = n4297_o;
  assign bus_en_flags_o = n4300_o;
  assign bus_write_sts_o = n4303_o;
  assign dm_write_dmem_addr_o = n4305_o;
  assign dm_write_dmem_o = n4577_o;
  assign dm_read_dmem_o = n4307_o;
  assign p1_write_p1_o = n4310_o;
  assign p1_read_p1_o = n4313_o;
  assign p2_write_p2_o = n4316_o;
  assign p2_write_exp_o = n4319_o;
  assign p2_read_p2_o = n4322_o;
  assign p2_read_exp_o = n4325_o;
  assign pm_write_pcl_o = n4328_o;
  assign pm_read_pcl_o = n4331_o;
  assign pm_write_pch_o = n4334_o;
  assign pm_read_pch_o = n4337_o;
  assign pm_read_pmem_o = n2110_o;
  assign psw_read_psw_o = n4340_o;
  assign psw_read_sp_o = n4343_o;
  assign psw_write_psw_o = n4346_o;
  assign psw_write_sp_o = n4349_o;
  assign alu_op_o = n4353_o;
  assign alu_use_carry_o = n4356_o;
  assign alu_da_high_o = n4359_o;
  assign alu_accu_low_o = n4362_o;
  assign alu_p06_temp_reg_o = n4365_o;
  assign alu_p60_temp_reg_o = n4368_o;
  assign bus_output_pcl_o = n2113_o;
  assign bus_bidir_bus_o = n4372_o;
  assign clk_multi_cycle_o = opc_multi_cycle_s;
  assign clk_assert_psen_o = n2116_o;
  assign clk_assert_prog_o = n4377_o;
  assign clk_assert_rd_o = n4381_o;
  assign clk_assert_wr_o = n4384_o;
  assign cnd_compute_take_o = n4387_o;
  assign cnd_branch_cond_o = n4397_o;
  assign cnd_comp_value_o = n4592_o;
  assign cnd_f1_o = f1_q;
  assign cnd_tf_o = tf_s;
  assign dm_addr_type_o = n4403_o;
  assign p1_read_reg_o = n4406_o;
  assign p2_read_reg_o = n4409_o;
  assign p2_output_pch_o = n2119_o;
  assign pm_inc_pc_o = n4578_o;
  assign pm_write_pmem_addr_o = n4579_o;
  assign pm_addr_type_o = n4412_o;
  assign psw_special_data_o = n4415_o;
  assign psw_inc_stackp_o = n4418_o;
  assign psw_dec_stackp_o = n4421_o;
  assign psw_write_carry_o = n4424_o;
  assign psw_write_aux_carry_o = n4427_o;
  assign psw_write_f0_o = n4430_o;
  assign psw_write_bs_o = n4433_o;
  assign tim_read_timer_o = n4436_o;
  assign tim_write_timer_o = n4439_o;
  assign tim_start_t_o = n4442_o;
  assign tim_start_cnt_o = n4445_o;
  assign tim_stop_tcnt_o = n4448_o;
  /* decoder.vhd:187:10  */
  assign opc_multi_cycle_s = n2006_o; // (signal)
  /* decoder.vhd:188:10  */
  assign opc_read_bus_s = n2122_o; // (signal)
  /* decoder.vhd:189:10  */
  assign opc_inj_int_s = n2125_o; // (signal)
  /* decoder.vhd:190:10  */
  assign opc_opcode_q = n4582_q; // (signal)
  /* decoder.vhd:191:10  */
  assign opc_mnemonic_s = n2008_o; // (signal)
  /* decoder.vhd:192:10  */
  assign last_cycle_s = n2026_o; // (signal)
  /* decoder.vhd:195:10  */
  assign assert_psen_s = n4473_o; // (signal)
  /* decoder.vhd:198:10  */
  assign branch_taken_s = n4476_o; // (signal)
  /* decoder.vhd:199:10  */
  assign branch_taken_q = n4584_q; // (signal)
  /* decoder.vhd:200:10  */
  assign pm_inc_pc_s = n2128_o; // (signal)
  /* decoder.vhd:201:10  */
  assign pm_write_pmem_addr_s = n2131_o; // (signal)
  /* decoder.vhd:203:10  */
  assign add_inc_pc_s = n4479_o; // (signal)
  /* decoder.vhd:205:10  */
  assign add_write_pmem_addr_s = n4482_o; // (signal)
  /* decoder.vhd:208:10  */
  assign clear_f1_s = n4485_o; // (signal)
  /* decoder.vhd:209:10  */
  assign cpl_f1_s = n4488_o; // (signal)
  /* decoder.vhd:210:10  */
  assign f1_q = n4585_q; // (signal)
  /* decoder.vhd:212:10  */
  assign clear_mb_s = n4491_o; // (signal)
  /* decoder.vhd:213:10  */
  assign set_mb_s = n4494_o; // (signal)
  /* decoder.vhd:214:10  */
  assign mb_q = n4587_q; // (signal)
  /* decoder.vhd:217:10  */
  assign ent0_clk_s = n4497_o; // (signal)
  /* decoder.vhd:218:10  */
  assign t0_dir_q = n4589_q; // (signal)
  /* decoder.vhd:220:10  */
  assign data_s = n4499_o; // (signal)
  /* decoder.vhd:221:10  */
  assign read_dec_s = n4500_o; // (signal)
  /* decoder.vhd:223:10  */
  assign tf_s = int_b_n2010; // (signal)
  /* decoder.vhd:225:10  */
  assign bus_read_bus_s = n2134_o; // (signal)
  /* decoder.vhd:226:10  */
  assign add_read_bus_s = n4502_o; // (signal)
  /* decoder.vhd:228:10  */
  assign dm_write_dmem_s = n4505_o; // (signal)
  /* decoder.vhd:230:10  */
  assign p2_output_exp_s = n4508_o; // (signal)
  /* decoder.vhd:232:10  */
  assign movx_first_cycle_s = n4511_o; // (signal)
  /* decoder.vhd:235:10  */
  assign jtf_executed_s = n4514_o; // (signal)
  /* decoder.vhd:236:10  */
  assign en_tcnti_s = n4517_o; // (signal)
  /* decoder.vhd:237:10  */
  assign dis_tcnti_s = n4520_o; // (signal)
  /* decoder.vhd:238:10  */
  assign en_i_s = n4523_o; // (signal)
  /* decoder.vhd:239:10  */
  assign dis_i_s = n4526_o; // (signal)
  /* decoder.vhd:240:10  */
  assign tim_int_s = int_b_n2012; // (signal)
  /* decoder.vhd:241:10  */
  assign retr_executed_s = n4529_o; // (signal)
  /* decoder.vhd:242:10  */
  assign int_executed_s = n4532_o; // (signal)
  /* decoder.vhd:243:10  */
  assign int_pending_s = int_b_n2013; // (signal)
  /* decoder.vhd:244:10  */
  assign int_in_progress_s = int_b_n2014; // (signal)
  /* decoder.vhd:247:10  */
  assign mnemonic_rec_s = n1986_o; // (signal)
  /* decoder.vhd:248:10  */
  assign mnemonic_q = n4591_q; // (signal)
  /* decoder_pack-p.vhd:553:7  */
  assign n1240_o = opc_opcode_q == 8'b11100101;
  /* decoder_pack-p.vhd:553:23  */
  assign n1242_o = opc_opcode_q == 8'b11110101;
  /* decoder_pack-p.vhd:553:23  */
  assign n1243_o = n1240_o | n1242_o;
  /* decoder_pack-p.vhd:558:7  */
  assign n1245_o = opc_opcode_q == 8'b10010000;
  assign n1246_o = {n1245_o, n1243_o};
  /* decoder_pack-p.vhd:551:5  */
  always @*
    case (n1246_o)
      2'b10: n1250_o = 6'b111111;
      2'b01: n1250_o = 6'b111110;
      default: n1250_o = 6'b000000;
    endcase
  /* decoder_pack-p.vhd:566:19  */
  assign n1253_o = n1250_o == 6'b000000;
  /* decoder_pack-p.vhd:491:7  */
  assign n1263_o = opc_opcode_q == 8'b10011001;
  /* decoder_pack-p.vhd:491:23  */
  assign n1265_o = opc_opcode_q == 8'b10011010;
  /* decoder_pack-p.vhd:491:23  */
  assign n1266_o = n1263_o | n1265_o;
  /* decoder_pack-p.vhd:496:7  */
  assign n1268_o = opc_opcode_q == 8'b00100010;
  /* decoder_pack-p.vhd:500:7  */
  assign n1270_o = opc_opcode_q == 8'b11010110;
  /* decoder_pack-p.vhd:505:7  */
  assign n1272_o = opc_opcode_q == 8'b10000110;
  /* decoder_pack-p.vhd:510:7  */
  assign n1274_o = opc_opcode_q == 8'b10001001;
  /* decoder_pack-p.vhd:510:23  */
  assign n1276_o = opc_opcode_q == 8'b10001010;
  /* decoder_pack-p.vhd:510:23  */
  assign n1277_o = n1274_o | n1276_o;
  /* decoder_pack-p.vhd:515:7  */
  assign n1279_o = opc_opcode_q == 8'b00000010;
  /* decoder_pack-p.vhd:519:7  */
  assign n1281_o = opc_opcode_q == 8'b00111001;
  /* decoder_pack-p.vhd:519:23  */
  assign n1283_o = opc_opcode_q == 8'b00111010;
  /* decoder_pack-p.vhd:519:23  */
  assign n1284_o = n1281_o | n1283_o;
  assign n1285_o = {n1284_o, n1279_o, n1277_o, n1272_o, n1270_o, n1268_o, n1266_o};
  /* decoder_pack-p.vhd:489:5  */
  always @*
    case (n1285_o)
      7'b1000000: n1294_o = 6'b101110;
      7'b0100000: n1294_o = 6'b111011;
      7'b0010000: n1294_o = 6'b101100;
      7'b0001000: n1294_o = 6'b111101;
      7'b0000100: n1294_o = 6'b111100;
      7'b0000010: n1294_o = 6'b111010;
      7'b0000001: n1294_o = 6'b000101;
      default: n1294_o = 6'b000000;
    endcase
  /* decoder_pack-p.vhd:489:5  */
  always @*
    case (n1285_o)
      7'b1000000: n1302_o = 1'b1;
      7'b0100000: n1302_o = 1'b0;
      7'b0010000: n1302_o = 1'b1;
      7'b0001000: n1302_o = 1'b1;
      7'b0000100: n1302_o = 1'b1;
      7'b0000010: n1302_o = 1'b0;
      7'b0000001: n1302_o = 1'b1;
      default: n1302_o = 1'b0;
    endcase
  /* decoder_pack-p.vhd:528:19  */
  assign n1305_o = n1294_o == 6'b000000;
  /* decoder_pack-p.vhd:123:7  */
  assign n1315_o = opc_opcode_q == 8'b01101000;
  /* decoder_pack-p.vhd:123:23  */
  assign n1317_o = opc_opcode_q == 8'b01101001;
  /* decoder_pack-p.vhd:123:23  */
  assign n1318_o = n1315_o | n1317_o;
  /* decoder_pack-p.vhd:123:36  */
  assign n1320_o = opc_opcode_q == 8'b01101010;
  /* decoder_pack-p.vhd:123:36  */
  assign n1321_o = n1318_o | n1320_o;
  /* decoder_pack-p.vhd:123:49  */
  assign n1323_o = opc_opcode_q == 8'b01101011;
  /* decoder_pack-p.vhd:123:49  */
  assign n1324_o = n1321_o | n1323_o;
  /* decoder_pack-p.vhd:123:62  */
  assign n1326_o = opc_opcode_q == 8'b01101100;
  /* decoder_pack-p.vhd:123:62  */
  assign n1327_o = n1324_o | n1326_o;
  /* decoder_pack-p.vhd:124:23  */
  assign n1329_o = opc_opcode_q == 8'b01101101;
  /* decoder_pack-p.vhd:124:23  */
  assign n1330_o = n1327_o | n1329_o;
  /* decoder_pack-p.vhd:124:36  */
  assign n1332_o = opc_opcode_q == 8'b01101110;
  /* decoder_pack-p.vhd:124:36  */
  assign n1333_o = n1330_o | n1332_o;
  /* decoder_pack-p.vhd:124:49  */
  assign n1335_o = opc_opcode_q == 8'b01101111;
  /* decoder_pack-p.vhd:124:49  */
  assign n1336_o = n1333_o | n1335_o;
  /* decoder_pack-p.vhd:124:62  */
  assign n1338_o = opc_opcode_q == 8'b01100000;
  /* decoder_pack-p.vhd:124:62  */
  assign n1339_o = n1336_o | n1338_o;
  /* decoder_pack-p.vhd:125:23  */
  assign n1341_o = opc_opcode_q == 8'b01100001;
  /* decoder_pack-p.vhd:125:23  */
  assign n1342_o = n1339_o | n1341_o;
  /* decoder_pack-p.vhd:125:36  */
  assign n1344_o = opc_opcode_q == 8'b01111000;
  /* decoder_pack-p.vhd:125:36  */
  assign n1345_o = n1342_o | n1344_o;
  /* decoder_pack-p.vhd:126:23  */
  assign n1347_o = opc_opcode_q == 8'b01111001;
  /* decoder_pack-p.vhd:126:23  */
  assign n1348_o = n1345_o | n1347_o;
  /* decoder_pack-p.vhd:126:36  */
  assign n1350_o = opc_opcode_q == 8'b01111010;
  /* decoder_pack-p.vhd:126:36  */
  assign n1351_o = n1348_o | n1350_o;
  /* decoder_pack-p.vhd:126:49  */
  assign n1353_o = opc_opcode_q == 8'b01111011;
  /* decoder_pack-p.vhd:126:49  */
  assign n1354_o = n1351_o | n1353_o;
  /* decoder_pack-p.vhd:126:62  */
  assign n1356_o = opc_opcode_q == 8'b01111100;
  /* decoder_pack-p.vhd:126:62  */
  assign n1357_o = n1354_o | n1356_o;
  /* decoder_pack-p.vhd:127:23  */
  assign n1359_o = opc_opcode_q == 8'b01111101;
  /* decoder_pack-p.vhd:127:23  */
  assign n1360_o = n1357_o | n1359_o;
  /* decoder_pack-p.vhd:127:36  */
  assign n1362_o = opc_opcode_q == 8'b01111110;
  /* decoder_pack-p.vhd:127:36  */
  assign n1363_o = n1360_o | n1362_o;
  /* decoder_pack-p.vhd:127:49  */
  assign n1365_o = opc_opcode_q == 8'b01111111;
  /* decoder_pack-p.vhd:127:49  */
  assign n1366_o = n1363_o | n1365_o;
  /* decoder_pack-p.vhd:127:62  */
  assign n1368_o = opc_opcode_q == 8'b01110000;
  /* decoder_pack-p.vhd:127:62  */
  assign n1369_o = n1366_o | n1368_o;
  /* decoder_pack-p.vhd:128:23  */
  assign n1371_o = opc_opcode_q == 8'b01110001;
  /* decoder_pack-p.vhd:128:23  */
  assign n1372_o = n1369_o | n1371_o;
  /* decoder_pack-p.vhd:132:7  */
  assign n1374_o = opc_opcode_q == 8'b00000011;
  /* decoder_pack-p.vhd:132:23  */
  assign n1376_o = opc_opcode_q == 8'b00010011;
  /* decoder_pack-p.vhd:132:23  */
  assign n1377_o = n1374_o | n1376_o;
  /* decoder_pack-p.vhd:138:7  */
  assign n1379_o = opc_opcode_q == 8'b01011000;
  /* decoder_pack-p.vhd:138:23  */
  assign n1381_o = opc_opcode_q == 8'b01011001;
  /* decoder_pack-p.vhd:138:23  */
  assign n1382_o = n1379_o | n1381_o;
  /* decoder_pack-p.vhd:138:36  */
  assign n1384_o = opc_opcode_q == 8'b01011010;
  /* decoder_pack-p.vhd:138:36  */
  assign n1385_o = n1382_o | n1384_o;
  /* decoder_pack-p.vhd:138:49  */
  assign n1387_o = opc_opcode_q == 8'b01011011;
  /* decoder_pack-p.vhd:138:49  */
  assign n1388_o = n1385_o | n1387_o;
  /* decoder_pack-p.vhd:138:62  */
  assign n1390_o = opc_opcode_q == 8'b01011100;
  /* decoder_pack-p.vhd:138:62  */
  assign n1391_o = n1388_o | n1390_o;
  /* decoder_pack-p.vhd:139:23  */
  assign n1393_o = opc_opcode_q == 8'b01011101;
  /* decoder_pack-p.vhd:139:23  */
  assign n1394_o = n1391_o | n1393_o;
  /* decoder_pack-p.vhd:139:36  */
  assign n1396_o = opc_opcode_q == 8'b01011110;
  /* decoder_pack-p.vhd:139:36  */
  assign n1397_o = n1394_o | n1396_o;
  /* decoder_pack-p.vhd:139:49  */
  assign n1399_o = opc_opcode_q == 8'b01011111;
  /* decoder_pack-p.vhd:139:49  */
  assign n1400_o = n1397_o | n1399_o;
  /* decoder_pack-p.vhd:139:62  */
  assign n1402_o = opc_opcode_q == 8'b01010000;
  /* decoder_pack-p.vhd:139:62  */
  assign n1403_o = n1400_o | n1402_o;
  /* decoder_pack-p.vhd:140:23  */
  assign n1405_o = opc_opcode_q == 8'b01010001;
  /* decoder_pack-p.vhd:140:23  */
  assign n1406_o = n1403_o | n1405_o;
  /* decoder_pack-p.vhd:144:7  */
  assign n1408_o = opc_opcode_q == 8'b01010011;
  /* decoder_pack-p.vhd:149:7  */
  assign n1410_o = opc_opcode_q == 8'b00010100;
  /* decoder_pack-p.vhd:149:23  */
  assign n1412_o = opc_opcode_q == 8'b00110100;
  /* decoder_pack-p.vhd:149:23  */
  assign n1413_o = n1410_o | n1412_o;
  /* decoder_pack-p.vhd:149:36  */
  assign n1415_o = opc_opcode_q == 8'b01010100;
  /* decoder_pack-p.vhd:149:36  */
  assign n1416_o = n1413_o | n1415_o;
  /* decoder_pack-p.vhd:149:49  */
  assign n1418_o = opc_opcode_q == 8'b01110100;
  /* decoder_pack-p.vhd:149:49  */
  assign n1419_o = n1416_o | n1418_o;
  /* decoder_pack-p.vhd:149:62  */
  assign n1421_o = opc_opcode_q == 8'b10010100;
  /* decoder_pack-p.vhd:149:62  */
  assign n1422_o = n1419_o | n1421_o;
  /* decoder_pack-p.vhd:150:23  */
  assign n1424_o = opc_opcode_q == 8'b10110100;
  /* decoder_pack-p.vhd:150:23  */
  assign n1425_o = n1422_o | n1424_o;
  /* decoder_pack-p.vhd:150:36  */
  assign n1427_o = opc_opcode_q == 8'b11010100;
  /* decoder_pack-p.vhd:150:36  */
  assign n1428_o = n1425_o | n1427_o;
  /* decoder_pack-p.vhd:150:49  */
  assign n1430_o = opc_opcode_q == 8'b11110100;
  /* decoder_pack-p.vhd:150:49  */
  assign n1431_o = n1428_o | n1430_o;
  /* decoder_pack-p.vhd:155:7  */
  assign n1433_o = opc_opcode_q == 8'b00100111;
  /* decoder_pack-p.vhd:159:7  */
  assign n1435_o = opc_opcode_q == 8'b10010111;
  /* decoder_pack-p.vhd:163:7  */
  assign n1437_o = opc_opcode_q == 8'b10000101;
  /* decoder_pack-p.vhd:163:23  */
  assign n1439_o = opc_opcode_q == 8'b10100101;
  /* decoder_pack-p.vhd:163:23  */
  assign n1440_o = n1437_o | n1439_o;
  /* decoder_pack-p.vhd:168:7  */
  assign n1442_o = opc_opcode_q == 8'b00110111;
  /* decoder_pack-p.vhd:172:7  */
  assign n1444_o = opc_opcode_q == 8'b10100111;
  /* decoder_pack-p.vhd:176:7  */
  assign n1446_o = opc_opcode_q == 8'b10010101;
  /* decoder_pack-p.vhd:176:23  */
  assign n1448_o = opc_opcode_q == 8'b10110101;
  /* decoder_pack-p.vhd:176:23  */
  assign n1449_o = n1446_o | n1448_o;
  /* decoder_pack-p.vhd:181:7  */
  assign n1451_o = opc_opcode_q == 8'b01010111;
  /* decoder_pack-p.vhd:185:7  */
  assign n1453_o = opc_opcode_q == 8'b11001000;
  /* decoder_pack-p.vhd:185:23  */
  assign n1455_o = opc_opcode_q == 8'b11001001;
  /* decoder_pack-p.vhd:185:23  */
  assign n1456_o = n1453_o | n1455_o;
  /* decoder_pack-p.vhd:185:36  */
  assign n1458_o = opc_opcode_q == 8'b11001010;
  /* decoder_pack-p.vhd:185:36  */
  assign n1459_o = n1456_o | n1458_o;
  /* decoder_pack-p.vhd:185:49  */
  assign n1461_o = opc_opcode_q == 8'b11001011;
  /* decoder_pack-p.vhd:185:49  */
  assign n1462_o = n1459_o | n1461_o;
  /* decoder_pack-p.vhd:185:62  */
  assign n1464_o = opc_opcode_q == 8'b11001100;
  /* decoder_pack-p.vhd:185:62  */
  assign n1465_o = n1462_o | n1464_o;
  /* decoder_pack-p.vhd:186:23  */
  assign n1467_o = opc_opcode_q == 8'b11001101;
  /* decoder_pack-p.vhd:186:23  */
  assign n1468_o = n1465_o | n1467_o;
  /* decoder_pack-p.vhd:186:36  */
  assign n1470_o = opc_opcode_q == 8'b11001110;
  /* decoder_pack-p.vhd:186:36  */
  assign n1471_o = n1468_o | n1470_o;
  /* decoder_pack-p.vhd:186:49  */
  assign n1473_o = opc_opcode_q == 8'b11001111;
  /* decoder_pack-p.vhd:186:49  */
  assign n1474_o = n1471_o | n1473_o;
  /* decoder_pack-p.vhd:186:62  */
  assign n1476_o = opc_opcode_q == 8'b00000111;
  /* decoder_pack-p.vhd:186:62  */
  assign n1477_o = n1474_o | n1476_o;
  /* decoder_pack-p.vhd:191:7  */
  assign n1479_o = opc_opcode_q == 8'b00010101;
  /* decoder_pack-p.vhd:191:23  */
  assign n1481_o = opc_opcode_q == 8'b00000101;
  /* decoder_pack-p.vhd:191:23  */
  assign n1482_o = n1479_o | n1481_o;
  /* decoder_pack-p.vhd:196:7  */
  assign n1484_o = opc_opcode_q == 8'b00110101;
  /* decoder_pack-p.vhd:196:23  */
  assign n1486_o = opc_opcode_q == 8'b00100101;
  /* decoder_pack-p.vhd:196:23  */
  assign n1487_o = n1484_o | n1486_o;
  /* decoder_pack-p.vhd:201:7  */
  assign n1489_o = opc_opcode_q == 8'b11101000;
  /* decoder_pack-p.vhd:201:23  */
  assign n1491_o = opc_opcode_q == 8'b11101001;
  /* decoder_pack-p.vhd:201:23  */
  assign n1492_o = n1489_o | n1491_o;
  /* decoder_pack-p.vhd:201:36  */
  assign n1494_o = opc_opcode_q == 8'b11101010;
  /* decoder_pack-p.vhd:201:36  */
  assign n1495_o = n1492_o | n1494_o;
  /* decoder_pack-p.vhd:201:49  */
  assign n1497_o = opc_opcode_q == 8'b11101011;
  /* decoder_pack-p.vhd:201:49  */
  assign n1498_o = n1495_o | n1497_o;
  /* decoder_pack-p.vhd:201:62  */
  assign n1500_o = opc_opcode_q == 8'b11101100;
  /* decoder_pack-p.vhd:201:62  */
  assign n1501_o = n1498_o | n1500_o;
  /* decoder_pack-p.vhd:202:23  */
  assign n1503_o = opc_opcode_q == 8'b11101101;
  /* decoder_pack-p.vhd:202:23  */
  assign n1504_o = n1501_o | n1503_o;
  /* decoder_pack-p.vhd:202:36  */
  assign n1506_o = opc_opcode_q == 8'b11101110;
  /* decoder_pack-p.vhd:202:36  */
  assign n1507_o = n1504_o | n1506_o;
  /* decoder_pack-p.vhd:202:49  */
  assign n1509_o = opc_opcode_q == 8'b11101111;
  /* decoder_pack-p.vhd:202:49  */
  assign n1510_o = n1507_o | n1509_o;
  /* decoder_pack-p.vhd:207:7  */
  assign n1512_o = opc_opcode_q == 8'b00001001;
  /* decoder_pack-p.vhd:207:23  */
  assign n1514_o = opc_opcode_q == 8'b00001010;
  /* decoder_pack-p.vhd:207:23  */
  assign n1515_o = n1512_o | n1514_o;
  /* decoder_pack-p.vhd:212:7  */
  assign n1517_o = opc_opcode_q == 8'b00010111;
  /* decoder_pack-p.vhd:212:23  */
  assign n1519_o = opc_opcode_q == 8'b00011000;
  /* decoder_pack-p.vhd:212:23  */
  assign n1520_o = n1517_o | n1519_o;
  /* decoder_pack-p.vhd:213:23  */
  assign n1522_o = opc_opcode_q == 8'b00011001;
  /* decoder_pack-p.vhd:213:23  */
  assign n1523_o = n1520_o | n1522_o;
  /* decoder_pack-p.vhd:213:36  */
  assign n1525_o = opc_opcode_q == 8'b00011010;
  /* decoder_pack-p.vhd:213:36  */
  assign n1526_o = n1523_o | n1525_o;
  /* decoder_pack-p.vhd:213:49  */
  assign n1528_o = opc_opcode_q == 8'b00011011;
  /* decoder_pack-p.vhd:213:49  */
  assign n1529_o = n1526_o | n1528_o;
  /* decoder_pack-p.vhd:213:62  */
  assign n1531_o = opc_opcode_q == 8'b00011100;
  /* decoder_pack-p.vhd:213:62  */
  assign n1532_o = n1529_o | n1531_o;
  /* decoder_pack-p.vhd:214:23  */
  assign n1534_o = opc_opcode_q == 8'b00011101;
  /* decoder_pack-p.vhd:214:23  */
  assign n1535_o = n1532_o | n1534_o;
  /* decoder_pack-p.vhd:214:36  */
  assign n1537_o = opc_opcode_q == 8'b00011110;
  /* decoder_pack-p.vhd:214:36  */
  assign n1538_o = n1535_o | n1537_o;
  /* decoder_pack-p.vhd:214:49  */
  assign n1540_o = opc_opcode_q == 8'b00011111;
  /* decoder_pack-p.vhd:214:49  */
  assign n1541_o = n1538_o | n1540_o;
  /* decoder_pack-p.vhd:214:62  */
  assign n1543_o = opc_opcode_q == 8'b00010000;
  /* decoder_pack-p.vhd:214:62  */
  assign n1544_o = n1541_o | n1543_o;
  /* decoder_pack-p.vhd:215:23  */
  assign n1546_o = opc_opcode_q == 8'b00010001;
  /* decoder_pack-p.vhd:215:23  */
  assign n1547_o = n1544_o | n1546_o;
  /* decoder_pack-p.vhd:219:7  */
  assign n1549_o = opc_opcode_q == 8'b00010010;
  /* decoder_pack-p.vhd:219:23  */
  assign n1551_o = opc_opcode_q == 8'b00110010;
  /* decoder_pack-p.vhd:219:23  */
  assign n1552_o = n1549_o | n1551_o;
  /* decoder_pack-p.vhd:219:36  */
  assign n1554_o = opc_opcode_q == 8'b01010010;
  /* decoder_pack-p.vhd:219:36  */
  assign n1555_o = n1552_o | n1554_o;
  /* decoder_pack-p.vhd:219:49  */
  assign n1557_o = opc_opcode_q == 8'b01110010;
  /* decoder_pack-p.vhd:219:49  */
  assign n1558_o = n1555_o | n1557_o;
  /* decoder_pack-p.vhd:219:62  */
  assign n1560_o = opc_opcode_q == 8'b10010010;
  /* decoder_pack-p.vhd:219:62  */
  assign n1561_o = n1558_o | n1560_o;
  /* decoder_pack-p.vhd:220:23  */
  assign n1563_o = opc_opcode_q == 8'b10110010;
  /* decoder_pack-p.vhd:220:23  */
  assign n1564_o = n1561_o | n1563_o;
  /* decoder_pack-p.vhd:220:36  */
  assign n1566_o = opc_opcode_q == 8'b11010010;
  /* decoder_pack-p.vhd:220:36  */
  assign n1567_o = n1564_o | n1566_o;
  /* decoder_pack-p.vhd:220:49  */
  assign n1569_o = opc_opcode_q == 8'b11110010;
  /* decoder_pack-p.vhd:220:49  */
  assign n1570_o = n1567_o | n1569_o;
  /* decoder_pack-p.vhd:225:7  */
  assign n1572_o = opc_opcode_q == 8'b11110110;
  /* decoder_pack-p.vhd:225:23  */
  assign n1574_o = opc_opcode_q == 8'b11100110;
  /* decoder_pack-p.vhd:225:23  */
  assign n1575_o = n1572_o | n1574_o;
  /* decoder_pack-p.vhd:231:7  */
  assign n1577_o = opc_opcode_q == 8'b10110110;
  /* decoder_pack-p.vhd:231:23  */
  assign n1579_o = opc_opcode_q == 8'b01110110;
  /* decoder_pack-p.vhd:231:23  */
  assign n1580_o = n1577_o | n1579_o;
  /* decoder_pack-p.vhd:237:7  */
  assign n1582_o = opc_opcode_q == 8'b00000100;
  /* decoder_pack-p.vhd:237:23  */
  assign n1584_o = opc_opcode_q == 8'b00100100;
  /* decoder_pack-p.vhd:237:23  */
  assign n1585_o = n1582_o | n1584_o;
  /* decoder_pack-p.vhd:237:36  */
  assign n1587_o = opc_opcode_q == 8'b01000100;
  /* decoder_pack-p.vhd:237:36  */
  assign n1588_o = n1585_o | n1587_o;
  /* decoder_pack-p.vhd:237:49  */
  assign n1590_o = opc_opcode_q == 8'b01100100;
  /* decoder_pack-p.vhd:237:49  */
  assign n1591_o = n1588_o | n1590_o;
  /* decoder_pack-p.vhd:237:62  */
  assign n1593_o = opc_opcode_q == 8'b10000100;
  /* decoder_pack-p.vhd:237:62  */
  assign n1594_o = n1591_o | n1593_o;
  /* decoder_pack-p.vhd:238:23  */
  assign n1596_o = opc_opcode_q == 8'b10100100;
  /* decoder_pack-p.vhd:238:23  */
  assign n1597_o = n1594_o | n1596_o;
  /* decoder_pack-p.vhd:238:36  */
  assign n1599_o = opc_opcode_q == 8'b11000100;
  /* decoder_pack-p.vhd:238:36  */
  assign n1600_o = n1597_o | n1599_o;
  /* decoder_pack-p.vhd:238:49  */
  assign n1602_o = opc_opcode_q == 8'b11100100;
  /* decoder_pack-p.vhd:238:49  */
  assign n1603_o = n1600_o | n1602_o;
  /* decoder_pack-p.vhd:243:7  */
  assign n1605_o = opc_opcode_q == 8'b10110011;
  /* decoder_pack-p.vhd:248:7  */
  assign n1607_o = opc_opcode_q == 8'b00100110;
  /* decoder_pack-p.vhd:248:23  */
  assign n1609_o = opc_opcode_q == 8'b01000110;
  /* decoder_pack-p.vhd:248:23  */
  assign n1610_o = n1607_o | n1609_o;
  /* decoder_pack-p.vhd:249:23  */
  assign n1612_o = opc_opcode_q == 8'b00110110;
  /* decoder_pack-p.vhd:249:23  */
  assign n1613_o = n1610_o | n1612_o;
  /* decoder_pack-p.vhd:250:23  */
  assign n1615_o = opc_opcode_q == 8'b01010110;
  /* decoder_pack-p.vhd:250:23  */
  assign n1616_o = n1613_o | n1615_o;
  /* decoder_pack-p.vhd:256:7  */
  assign n1618_o = opc_opcode_q == 8'b00010110;
  /* decoder_pack-p.vhd:261:7  */
  assign n1620_o = opc_opcode_q == 8'b10010110;
  /* decoder_pack-p.vhd:261:23  */
  assign n1622_o = opc_opcode_q == 8'b11000110;
  /* decoder_pack-p.vhd:261:23  */
  assign n1623_o = n1620_o | n1622_o;
  /* decoder_pack-p.vhd:267:7  */
  assign n1625_o = opc_opcode_q == 8'b00100011;
  /* decoder_pack-p.vhd:272:7  */
  assign n1627_o = opc_opcode_q == 8'b11000111;
  /* decoder_pack-p.vhd:276:7  */
  assign n1629_o = opc_opcode_q == 8'b11111000;
  /* decoder_pack-p.vhd:276:23  */
  assign n1631_o = opc_opcode_q == 8'b11111001;
  /* decoder_pack-p.vhd:276:23  */
  assign n1632_o = n1629_o | n1631_o;
  /* decoder_pack-p.vhd:276:36  */
  assign n1634_o = opc_opcode_q == 8'b11111010;
  /* decoder_pack-p.vhd:276:36  */
  assign n1635_o = n1632_o | n1634_o;
  /* decoder_pack-p.vhd:276:49  */
  assign n1637_o = opc_opcode_q == 8'b11111011;
  /* decoder_pack-p.vhd:276:49  */
  assign n1638_o = n1635_o | n1637_o;
  /* decoder_pack-p.vhd:276:62  */
  assign n1640_o = opc_opcode_q == 8'b11111100;
  /* decoder_pack-p.vhd:276:62  */
  assign n1641_o = n1638_o | n1640_o;
  /* decoder_pack-p.vhd:277:23  */
  assign n1643_o = opc_opcode_q == 8'b11111101;
  /* decoder_pack-p.vhd:277:23  */
  assign n1644_o = n1641_o | n1643_o;
  /* decoder_pack-p.vhd:277:36  */
  assign n1646_o = opc_opcode_q == 8'b11111110;
  /* decoder_pack-p.vhd:277:36  */
  assign n1647_o = n1644_o | n1646_o;
  /* decoder_pack-p.vhd:277:49  */
  assign n1649_o = opc_opcode_q == 8'b11111111;
  /* decoder_pack-p.vhd:277:49  */
  assign n1650_o = n1647_o | n1649_o;
  /* decoder_pack-p.vhd:277:62  */
  assign n1652_o = opc_opcode_q == 8'b11110000;
  /* decoder_pack-p.vhd:277:62  */
  assign n1653_o = n1650_o | n1652_o;
  /* decoder_pack-p.vhd:278:23  */
  assign n1655_o = opc_opcode_q == 8'b11110001;
  /* decoder_pack-p.vhd:278:23  */
  assign n1656_o = n1653_o | n1655_o;
  /* decoder_pack-p.vhd:282:7  */
  assign n1658_o = opc_opcode_q == 8'b11010111;
  /* decoder_pack-p.vhd:286:7  */
  assign n1660_o = opc_opcode_q == 8'b10101000;
  /* decoder_pack-p.vhd:286:23  */
  assign n1662_o = opc_opcode_q == 8'b10101001;
  /* decoder_pack-p.vhd:286:23  */
  assign n1663_o = n1660_o | n1662_o;
  /* decoder_pack-p.vhd:286:36  */
  assign n1665_o = opc_opcode_q == 8'b10101010;
  /* decoder_pack-p.vhd:286:36  */
  assign n1666_o = n1663_o | n1665_o;
  /* decoder_pack-p.vhd:286:49  */
  assign n1668_o = opc_opcode_q == 8'b10101011;
  /* decoder_pack-p.vhd:286:49  */
  assign n1669_o = n1666_o | n1668_o;
  /* decoder_pack-p.vhd:286:62  */
  assign n1671_o = opc_opcode_q == 8'b10101100;
  /* decoder_pack-p.vhd:286:62  */
  assign n1672_o = n1669_o | n1671_o;
  /* decoder_pack-p.vhd:287:23  */
  assign n1674_o = opc_opcode_q == 8'b10101101;
  /* decoder_pack-p.vhd:287:23  */
  assign n1675_o = n1672_o | n1674_o;
  /* decoder_pack-p.vhd:287:36  */
  assign n1677_o = opc_opcode_q == 8'b10101110;
  /* decoder_pack-p.vhd:287:36  */
  assign n1678_o = n1675_o | n1677_o;
  /* decoder_pack-p.vhd:287:49  */
  assign n1680_o = opc_opcode_q == 8'b10101111;
  /* decoder_pack-p.vhd:287:49  */
  assign n1681_o = n1678_o | n1680_o;
  /* decoder_pack-p.vhd:287:62  */
  assign n1683_o = opc_opcode_q == 8'b10100000;
  /* decoder_pack-p.vhd:287:62  */
  assign n1684_o = n1681_o | n1683_o;
  /* decoder_pack-p.vhd:288:23  */
  assign n1686_o = opc_opcode_q == 8'b10100001;
  /* decoder_pack-p.vhd:288:23  */
  assign n1687_o = n1684_o | n1686_o;
  /* decoder_pack-p.vhd:292:7  */
  assign n1689_o = opc_opcode_q == 8'b10111000;
  /* decoder_pack-p.vhd:292:23  */
  assign n1691_o = opc_opcode_q == 8'b10111001;
  /* decoder_pack-p.vhd:292:23  */
  assign n1692_o = n1689_o | n1691_o;
  /* decoder_pack-p.vhd:292:36  */
  assign n1694_o = opc_opcode_q == 8'b10111010;
  /* decoder_pack-p.vhd:292:36  */
  assign n1695_o = n1692_o | n1694_o;
  /* decoder_pack-p.vhd:292:49  */
  assign n1697_o = opc_opcode_q == 8'b10111011;
  /* decoder_pack-p.vhd:292:49  */
  assign n1698_o = n1695_o | n1697_o;
  /* decoder_pack-p.vhd:292:62  */
  assign n1700_o = opc_opcode_q == 8'b10111100;
  /* decoder_pack-p.vhd:292:62  */
  assign n1701_o = n1698_o | n1700_o;
  /* decoder_pack-p.vhd:293:23  */
  assign n1703_o = opc_opcode_q == 8'b10111101;
  /* decoder_pack-p.vhd:293:23  */
  assign n1704_o = n1701_o | n1703_o;
  /* decoder_pack-p.vhd:293:36  */
  assign n1706_o = opc_opcode_q == 8'b10111110;
  /* decoder_pack-p.vhd:293:36  */
  assign n1707_o = n1704_o | n1706_o;
  /* decoder_pack-p.vhd:293:49  */
  assign n1709_o = opc_opcode_q == 8'b10111111;
  /* decoder_pack-p.vhd:293:49  */
  assign n1710_o = n1707_o | n1709_o;
  /* decoder_pack-p.vhd:293:62  */
  assign n1712_o = opc_opcode_q == 8'b10110000;
  /* decoder_pack-p.vhd:293:62  */
  assign n1713_o = n1710_o | n1712_o;
  /* decoder_pack-p.vhd:294:23  */
  assign n1715_o = opc_opcode_q == 8'b10110001;
  /* decoder_pack-p.vhd:294:23  */
  assign n1716_o = n1713_o | n1715_o;
  /* decoder_pack-p.vhd:299:7  */
  assign n1718_o = opc_opcode_q == 8'b01100010;
  /* decoder_pack-p.vhd:299:23  */
  assign n1720_o = opc_opcode_q == 8'b01000010;
  /* decoder_pack-p.vhd:299:23  */
  assign n1721_o = n1718_o | n1720_o;
  /* decoder_pack-p.vhd:304:7  */
  assign n1723_o = opc_opcode_q == 8'b00001100;
  /* decoder_pack-p.vhd:304:23  */
  assign n1725_o = opc_opcode_q == 8'b00001101;
  /* decoder_pack-p.vhd:304:23  */
  assign n1726_o = n1723_o | n1725_o;
  /* decoder_pack-p.vhd:304:36  */
  assign n1728_o = opc_opcode_q == 8'b00001110;
  /* decoder_pack-p.vhd:304:36  */
  assign n1729_o = n1726_o | n1728_o;
  /* decoder_pack-p.vhd:304:49  */
  assign n1731_o = opc_opcode_q == 8'b00001111;
  /* decoder_pack-p.vhd:304:49  */
  assign n1732_o = n1729_o | n1731_o;
  /* decoder_pack-p.vhd:309:7  */
  assign n1734_o = opc_opcode_q == 8'b10100011;
  /* decoder_pack-p.vhd:309:23  */
  assign n1736_o = opc_opcode_q == 8'b11100011;
  /* decoder_pack-p.vhd:309:23  */
  assign n1737_o = n1734_o | n1736_o;
  /* decoder_pack-p.vhd:315:7  */
  assign n1739_o = opc_opcode_q == 8'b00000000;
  /* decoder_pack-p.vhd:319:7  */
  assign n1741_o = opc_opcode_q == 8'b01001000;
  /* decoder_pack-p.vhd:319:23  */
  assign n1743_o = opc_opcode_q == 8'b01001001;
  /* decoder_pack-p.vhd:319:23  */
  assign n1744_o = n1741_o | n1743_o;
  /* decoder_pack-p.vhd:319:36  */
  assign n1746_o = opc_opcode_q == 8'b01001010;
  /* decoder_pack-p.vhd:319:36  */
  assign n1747_o = n1744_o | n1746_o;
  /* decoder_pack-p.vhd:319:49  */
  assign n1749_o = opc_opcode_q == 8'b01001011;
  /* decoder_pack-p.vhd:319:49  */
  assign n1750_o = n1747_o | n1749_o;
  /* decoder_pack-p.vhd:319:62  */
  assign n1752_o = opc_opcode_q == 8'b01001100;
  /* decoder_pack-p.vhd:319:62  */
  assign n1753_o = n1750_o | n1752_o;
  /* decoder_pack-p.vhd:320:23  */
  assign n1755_o = opc_opcode_q == 8'b01001101;
  /* decoder_pack-p.vhd:320:23  */
  assign n1756_o = n1753_o | n1755_o;
  /* decoder_pack-p.vhd:320:36  */
  assign n1758_o = opc_opcode_q == 8'b01001110;
  /* decoder_pack-p.vhd:320:36  */
  assign n1759_o = n1756_o | n1758_o;
  /* decoder_pack-p.vhd:320:49  */
  assign n1761_o = opc_opcode_q == 8'b01001111;
  /* decoder_pack-p.vhd:320:49  */
  assign n1762_o = n1759_o | n1761_o;
  /* decoder_pack-p.vhd:320:62  */
  assign n1764_o = opc_opcode_q == 8'b01000000;
  /* decoder_pack-p.vhd:320:62  */
  assign n1765_o = n1762_o | n1764_o;
  /* decoder_pack-p.vhd:321:23  */
  assign n1767_o = opc_opcode_q == 8'b01000001;
  /* decoder_pack-p.vhd:321:23  */
  assign n1768_o = n1765_o | n1767_o;
  /* decoder_pack-p.vhd:325:7  */
  assign n1770_o = opc_opcode_q == 8'b01000011;
  /* decoder_pack-p.vhd:330:7  */
  assign n1772_o = opc_opcode_q == 8'b00111100;
  /* decoder_pack-p.vhd:330:23  */
  assign n1774_o = opc_opcode_q == 8'b00111101;
  /* decoder_pack-p.vhd:330:23  */
  assign n1775_o = n1772_o | n1774_o;
  /* decoder_pack-p.vhd:330:36  */
  assign n1777_o = opc_opcode_q == 8'b00111110;
  /* decoder_pack-p.vhd:330:36  */
  assign n1778_o = n1775_o | n1777_o;
  /* decoder_pack-p.vhd:330:49  */
  assign n1780_o = opc_opcode_q == 8'b00111111;
  /* decoder_pack-p.vhd:330:49  */
  assign n1781_o = n1778_o | n1780_o;
  /* decoder_pack-p.vhd:330:62  */
  assign n1783_o = opc_opcode_q == 8'b10011100;
  /* decoder_pack-p.vhd:330:62  */
  assign n1784_o = n1781_o | n1783_o;
  /* decoder_pack-p.vhd:331:23  */
  assign n1786_o = opc_opcode_q == 8'b10011101;
  /* decoder_pack-p.vhd:331:23  */
  assign n1787_o = n1784_o | n1786_o;
  /* decoder_pack-p.vhd:331:36  */
  assign n1789_o = opc_opcode_q == 8'b10011110;
  /* decoder_pack-p.vhd:331:36  */
  assign n1790_o = n1787_o | n1789_o;
  /* decoder_pack-p.vhd:331:49  */
  assign n1792_o = opc_opcode_q == 8'b10011111;
  /* decoder_pack-p.vhd:331:49  */
  assign n1793_o = n1790_o | n1792_o;
  /* decoder_pack-p.vhd:331:62  */
  assign n1795_o = opc_opcode_q == 8'b10001100;
  /* decoder_pack-p.vhd:331:62  */
  assign n1796_o = n1793_o | n1795_o;
  /* decoder_pack-p.vhd:332:23  */
  assign n1798_o = opc_opcode_q == 8'b10001101;
  /* decoder_pack-p.vhd:332:23  */
  assign n1799_o = n1796_o | n1798_o;
  /* decoder_pack-p.vhd:332:36  */
  assign n1801_o = opc_opcode_q == 8'b10001110;
  /* decoder_pack-p.vhd:332:36  */
  assign n1802_o = n1799_o | n1801_o;
  /* decoder_pack-p.vhd:332:49  */
  assign n1804_o = opc_opcode_q == 8'b10001111;
  /* decoder_pack-p.vhd:332:49  */
  assign n1805_o = n1802_o | n1804_o;
  /* decoder_pack-p.vhd:337:7  */
  assign n1807_o = opc_opcode_q == 8'b10000011;
  /* decoder_pack-p.vhd:337:23  */
  assign n1809_o = opc_opcode_q == 8'b10010011;
  /* decoder_pack-p.vhd:337:23  */
  assign n1810_o = n1807_o | n1809_o;
  /* decoder_pack-p.vhd:343:7  */
  assign n1812_o = opc_opcode_q == 8'b11100111;
  /* decoder_pack-p.vhd:343:23  */
  assign n1814_o = opc_opcode_q == 8'b11110111;
  /* decoder_pack-p.vhd:343:23  */
  assign n1815_o = n1812_o | n1814_o;
  /* decoder_pack-p.vhd:348:7  */
  assign n1817_o = opc_opcode_q == 8'b01110111;
  /* decoder_pack-p.vhd:348:23  */
  assign n1819_o = opc_opcode_q == 8'b01100111;
  /* decoder_pack-p.vhd:348:23  */
  assign n1820_o = n1817_o | n1819_o;
  /* decoder_pack-p.vhd:353:7  */
  assign n1822_o = opc_opcode_q == 8'b11000101;
  /* decoder_pack-p.vhd:353:23  */
  assign n1824_o = opc_opcode_q == 8'b11010101;
  /* decoder_pack-p.vhd:353:23  */
  assign n1825_o = n1822_o | n1824_o;
  /* decoder_pack-p.vhd:358:7  */
  assign n1827_o = opc_opcode_q == 8'b01100101;
  /* decoder_pack-p.vhd:362:7  */
  assign n1829_o = opc_opcode_q == 8'b01000101;
  /* decoder_pack-p.vhd:362:23  */
  assign n1831_o = opc_opcode_q == 8'b01010101;
  /* decoder_pack-p.vhd:362:23  */
  assign n1832_o = n1829_o | n1831_o;
  /* decoder_pack-p.vhd:367:7  */
  assign n1834_o = opc_opcode_q == 8'b01000111;
  /* decoder_pack-p.vhd:371:7  */
  assign n1836_o = opc_opcode_q == 8'b00101000;
  /* decoder_pack-p.vhd:371:23  */
  assign n1838_o = opc_opcode_q == 8'b00101001;
  /* decoder_pack-p.vhd:371:23  */
  assign n1839_o = n1836_o | n1838_o;
  /* decoder_pack-p.vhd:371:36  */
  assign n1841_o = opc_opcode_q == 8'b00101010;
  /* decoder_pack-p.vhd:371:36  */
  assign n1842_o = n1839_o | n1841_o;
  /* decoder_pack-p.vhd:371:49  */
  assign n1844_o = opc_opcode_q == 8'b00101011;
  /* decoder_pack-p.vhd:371:49  */
  assign n1845_o = n1842_o | n1844_o;
  /* decoder_pack-p.vhd:371:62  */
  assign n1847_o = opc_opcode_q == 8'b00101100;
  /* decoder_pack-p.vhd:371:62  */
  assign n1848_o = n1845_o | n1847_o;
  /* decoder_pack-p.vhd:372:23  */
  assign n1850_o = opc_opcode_q == 8'b00101101;
  /* decoder_pack-p.vhd:372:23  */
  assign n1851_o = n1848_o | n1850_o;
  /* decoder_pack-p.vhd:372:36  */
  assign n1853_o = opc_opcode_q == 8'b00101110;
  /* decoder_pack-p.vhd:372:36  */
  assign n1854_o = n1851_o | n1853_o;
  /* decoder_pack-p.vhd:372:49  */
  assign n1856_o = opc_opcode_q == 8'b00101111;
  /* decoder_pack-p.vhd:372:49  */
  assign n1857_o = n1854_o | n1856_o;
  /* decoder_pack-p.vhd:372:62  */
  assign n1859_o = opc_opcode_q == 8'b00100000;
  /* decoder_pack-p.vhd:372:62  */
  assign n1860_o = n1857_o | n1859_o;
  /* decoder_pack-p.vhd:373:23  */
  assign n1862_o = opc_opcode_q == 8'b00100001;
  /* decoder_pack-p.vhd:373:23  */
  assign n1863_o = n1860_o | n1862_o;
  /* decoder_pack-p.vhd:373:36  */
  assign n1865_o = opc_opcode_q == 8'b00110000;
  /* decoder_pack-p.vhd:373:36  */
  assign n1866_o = n1863_o | n1865_o;
  /* decoder_pack-p.vhd:374:23  */
  assign n1868_o = opc_opcode_q == 8'b00110001;
  /* decoder_pack-p.vhd:374:23  */
  assign n1869_o = n1866_o | n1868_o;
  /* decoder_pack-p.vhd:378:7  */
  assign n1871_o = opc_opcode_q == 8'b11011000;
  /* decoder_pack-p.vhd:378:23  */
  assign n1873_o = opc_opcode_q == 8'b11011001;
  /* decoder_pack-p.vhd:378:23  */
  assign n1874_o = n1871_o | n1873_o;
  /* decoder_pack-p.vhd:378:36  */
  assign n1876_o = opc_opcode_q == 8'b11011010;
  /* decoder_pack-p.vhd:378:36  */
  assign n1877_o = n1874_o | n1876_o;
  /* decoder_pack-p.vhd:378:49  */
  assign n1879_o = opc_opcode_q == 8'b11011011;
  /* decoder_pack-p.vhd:378:49  */
  assign n1880_o = n1877_o | n1879_o;
  /* decoder_pack-p.vhd:378:62  */
  assign n1882_o = opc_opcode_q == 8'b11011100;
  /* decoder_pack-p.vhd:378:62  */
  assign n1883_o = n1880_o | n1882_o;
  /* decoder_pack-p.vhd:379:23  */
  assign n1885_o = opc_opcode_q == 8'b11011101;
  /* decoder_pack-p.vhd:379:23  */
  assign n1886_o = n1883_o | n1885_o;
  /* decoder_pack-p.vhd:379:36  */
  assign n1888_o = opc_opcode_q == 8'b11011110;
  /* decoder_pack-p.vhd:379:36  */
  assign n1889_o = n1886_o | n1888_o;
  /* decoder_pack-p.vhd:379:49  */
  assign n1891_o = opc_opcode_q == 8'b11011111;
  /* decoder_pack-p.vhd:379:49  */
  assign n1892_o = n1889_o | n1891_o;
  /* decoder_pack-p.vhd:379:62  */
  assign n1894_o = opc_opcode_q == 8'b11010000;
  /* decoder_pack-p.vhd:379:62  */
  assign n1895_o = n1892_o | n1894_o;
  /* decoder_pack-p.vhd:380:23  */
  assign n1897_o = opc_opcode_q == 8'b11010001;
  /* decoder_pack-p.vhd:380:23  */
  assign n1898_o = n1895_o | n1897_o;
  /* decoder_pack-p.vhd:384:7  */
  assign n1900_o = opc_opcode_q == 8'b11010011;
  assign n1901_o = {n1900_o, n1898_o, n1869_o, n1834_o, n1832_o, n1827_o, n1825_o, n1820_o, n1815_o, n1810_o, n1805_o, n1770_o, n1768_o, n1739_o, n1737_o, n1732_o, n1721_o, n1716_o, n1687_o, n1658_o, n1656_o, n1627_o, n1625_o, n1623_o, n1618_o, n1616_o, n1605_o, n1603_o, n1580_o, n1575_o, n1570_o, n1547_o, n1515_o, n1510_o, n1487_o, n1482_o, n1477_o, n1451_o, n1449_o, n1444_o, n1442_o, n1440_o, n1435_o, n1433_o, n1431_o, n1408_o, n1406_o, n1377_o, n1372_o};
  /* decoder_pack-p.vhd:121:5  */
  always @*
    case (n1901_o)
      49'b1000000000000000000000000000000000000000000000000: n1952_o = 6'b111001;
      49'b0100000000000000000000000000000000000000000000000: n1952_o = 6'b111000;
      49'b0010000000000000000000000000000000000000000000000: n1952_o = 6'b110111;
      49'b0001000000000000000000000000000000000000000000000: n1952_o = 6'b110110;
      49'b0000100000000000000000000000000000000000000000000: n1952_o = 6'b110101;
      49'b0000010000000000000000000000000000000000000000000: n1952_o = 6'b110100;
      49'b0000001000000000000000000000000000000000000000000: n1952_o = 6'b110011;
      49'b0000000100000000000000000000000000000000000000000: n1952_o = 6'b110001;
      49'b0000000010000000000000000000000000000000000000000: n1952_o = 6'b110000;
      49'b0000000001000000000000000000000000000000000000000: n1952_o = 6'b101111;
      49'b0000000000100000000000000000000000000000000000000: n1952_o = 6'b101101;
      49'b0000000000010000000000000000000000000000000000000: n1952_o = 6'b101011;
      49'b0000000000001000000000000000000000000000000000000: n1952_o = 6'b101010;
      49'b0000000000000100000000000000000000000000000000000: n1952_o = 6'b101001;
      49'b0000000000000010000000000000000000000000000000000: n1952_o = 6'b100111;
      49'b0000000000000001000000000000000000000000000000000: n1952_o = 6'b100110;
      49'b0000000000000000100000000000000000000000000000000: n1952_o = 6'b100101;
      49'b0000000000000000010000000000000000000000000000000: n1952_o = 6'b100100;
      49'b0000000000000000001000000000000000000000000000000: n1952_o = 6'b100011;
      49'b0000000000000000000100000000000000000000000000000: n1952_o = 6'b100010;
      49'b0000000000000000000010000000000000000000000000000: n1952_o = 6'b100001;
      49'b0000000000000000000001000000000000000000000000000: n1952_o = 6'b100000;
      49'b0000000000000000000000100000000000000000000000000: n1952_o = 6'b011111;
      49'b0000000000000000000000010000000000000000000000000: n1952_o = 6'b011110;
      49'b0000000000000000000000001000000000000000000000000: n1952_o = 6'b011101;
      49'b0000000000000000000000000100000000000000000000000: n1952_o = 6'b011100;
      49'b0000000000000000000000000010000000000000000000000: n1952_o = 6'b011010;
      49'b0000000000000000000000000001000000000000000000000: n1952_o = 6'b011001;
      49'b0000000000000000000000000000100000000000000000000: n1952_o = 6'b011000;
      49'b0000000000000000000000000000010000000000000000000: n1952_o = 6'b010111;
      49'b0000000000000000000000000000001000000000000000000: n1952_o = 6'b010110;
      49'b0000000000000000000000000000000100000000000000000: n1952_o = 6'b010100;
      49'b0000000000000000000000000000000010000000000000000: n1952_o = 6'b010011;
      49'b0000000000000000000000000000000001000000000000000: n1952_o = 6'b010001;
      49'b0000000000000000000000000000000000100000000000000: n1952_o = 6'b010000;
      49'b0000000000000000000000000000000000010000000000000: n1952_o = 6'b001111;
      49'b0000000000000000000000000000000000001000000000000: n1952_o = 6'b001110;
      49'b0000000000000000000000000000000000000100000000000: n1952_o = 6'b001101;
      49'b0000000000000000000000000000000000000010000000000: n1952_o = 6'b001100;
      49'b0000000000000000000000000000000000000001000000000: n1952_o = 6'b001011;
      49'b0000000000000000000000000000000000000000100000000: n1952_o = 6'b001010;
      49'b0000000000000000000000000000000000000000010000000: n1952_o = 6'b001001;
      49'b0000000000000000000000000000000000000000001000000: n1952_o = 6'b001000;
      49'b0000000000000000000000000000000000000000000100000: n1952_o = 6'b000111;
      49'b0000000000000000000000000000000000000000000010000: n1952_o = 6'b000110;
      49'b0000000000000000000000000000000000000000000001000: n1952_o = 6'b000100;
      49'b0000000000000000000000000000000000000000000000100: n1952_o = 6'b000011;
      49'b0000000000000000000000000000000000000000000000010: n1952_o = 6'b000010;
      49'b0000000000000000000000000000000000000000000000001: n1952_o = 6'b000001;
      default: n1952_o = 6'b101001;
    endcase
  /* decoder_pack-p.vhd:121:5  */
  always @*
    case (n1901_o)
      49'b1000000000000000000000000000000000000000000000000: n1976_o = 1'b1;
      49'b0100000000000000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0010000000000000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0001000000000000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000100000000000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000010000000000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000001000000000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000100000000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000010000000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000001000000000000000000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000100000000000000000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000010000000000000000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000001000000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000000000100000000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000000000010000000000000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000001000000000000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000100000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000000000000010000000000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000001000000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000000000000000100000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000000000000000010000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000000000000000001000000000000000000000000000: n1976_o = 1'b0;
      49'b0000000000000000000000100000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000010000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000001000000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000100000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000010000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000001000000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000000100000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000000010000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000000001000000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000000000100000000000000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000010000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000000000001000000000000000: n1976_o = 1'b1;
      49'b0000000000000000000000000000000000100000000000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000010000000000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000001000000000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000100000000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000010000000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000001000000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000000100000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000000010000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000000001000000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000000000100000: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000000000010000: n1976_o = 1'b1;
      49'b0000000000000000000000000000000000000000000001000: n1976_o = 1'b1;
      49'b0000000000000000000000000000000000000000000000100: n1976_o = 1'b0;
      49'b0000000000000000000000000000000000000000000000010: n1976_o = 1'b1;
      49'b0000000000000000000000000000000000000000000000001: n1976_o = 1'b0;
      default: n1976_o = 1'b0;
    endcase
  assign n1980_o = {n1976_o, n1952_o};
  assign n1981_o = {n1302_o, n1294_o};
  /* decoder_pack-p.vhd:528:5  */
  assign n1982_o = n1305_o ? n1980_o : n1981_o;
  assign n1985_o = {1'b0, n1250_o};
  /* decoder_pack-p.vhd:566:5  */
  assign n1986_o = n1253_o ? n1982_o : n1985_o;
  /* decoder.vhd:301:14  */
  assign n1989_o = ~res_i;
  /* decoder.vhd:313:40  */
  assign n1991_o = mnemonic_rec_s[5:0];
  /* decoder.vhd:310:9  */
  assign n1993_o = opc_inj_int_s ? 8'b00010100 : opc_opcode_q;
  /* decoder.vhd:310:9  */
  assign n1994_o = opc_inj_int_s ? mnemonic_q : n1991_o;
  /* decoder.vhd:308:9  */
  assign n1995_o = opc_read_bus_s ? data_i : n1993_o;
  /* decoder.vhd:308:9  */
  assign n1996_o = opc_read_bus_s ? mnemonic_q : n1994_o;
  /* decoder.vhd:322:39  */
  assign n2006_o = mnemonic_rec_s[6];
  /* decoder.vhd:324:24  */
  assign n2008_o = 1'b1 ? mnemonic_q : n2009_o;
  /* decoder.vhd:325:41  */
  assign n2009_o = mnemonic_rec_s[5:0];
  /* decoder.vhd:343:28  */
  assign int_b_n2010 = int_b_tf_o; // (signal)
  /* decoder.vhd:352:28  */
  assign int_b_n2012 = int_b_tim_int_o; // (signal)
  /* decoder.vhd:355:28  */
  assign int_b_n2013 = int_b_int_pending_o; // (signal)
  /* decoder.vhd:356:28  */
  assign int_b_n2014 = int_b_int_in_progress_o; // (signal)
  /* decoder.vhd:333:3  */
  t48_int int_b (
    .clk_i(clk_i),
    .res_i(res_i),
    .en_clk_i(en_clk_i),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_i),
    .clk_mstate_i(clk_mstate_i),
    .jtf_executed_i(jtf_executed_s),
    .tim_overflow_i(tim_overflow_i),
    .en_tcnti_i(en_tcnti_s),
    .dis_tcnti_i(dis_tcnti_s),
    .int_n_i(int_n_i),
    .ale_i(ale_i),
    .last_cycle_i(last_cycle_s),
    .en_i_i(en_i_s),
    .dis_i_i(dis_i_s),
    .retr_executed_i(retr_executed_s),
    .int_executed_i(int_executed_s),
    .tf_o(int_b_tf_o),
    .ext_int_o(),
    .tim_int_o(int_b_tim_int_o),
    .int_pending_o(int_b_int_pending_o),
    .int_in_progress_o(int_b_int_in_progress_o));
  /* decoder.vhd:359:19  */
  assign n2024_o = ~opc_multi_cycle_s;
  /* decoder.vhd:360:38  */
  assign n2025_o = opc_multi_cycle_s & clk_second_cycle_i;
  /* decoder.vhd:359:41  */
  assign n2026_o = n2024_o | n2025_o;
  /* decoder.vhd:393:26  */
  assign n2029_o = ~clk_second_cycle_i;
  /* decoder.vhd:394:46  */
  assign n2030_o = clk_second_cycle_i & assert_psen_s;
  /* decoder.vhd:393:49  */
  assign n2031_o = n2029_o | n2030_o;
  /* decoder.vhd:399:19  */
  assign n2032_o = ~ea_i;
  /* decoder.vhd:400:16  */
  assign n2033_o = ~int_pending_s;
  /* decoder.vhd:400:13  */
  assign n2036_o = n2033_o ? 1'b1 : 1'b0;
  /* decoder.vhd:405:16  */
  assign n2037_o = ~int_pending_s;
  /* decoder.vhd:405:13  */
  assign n2040_o = n2037_o ? 1'b1 : 1'b0;
  /* decoder.vhd:399:11  */
  assign n2042_o = n2032_o ? n2036_o : 1'b0;
  /* decoder.vhd:399:11  */
  assign n2045_o = n2032_o ? 1'b0 : 1'b1;
  /* decoder.vhd:399:11  */
  assign n2047_o = n2032_o ? 1'b0 : n2040_o;
  /* decoder.vhd:398:9  */
  assign n2049_o = n2031_o ? n2042_o : 1'b0;
  /* decoder.vhd:398:9  */
  assign n2051_o = n2031_o ? n2045_o : 1'b0;
  /* decoder.vhd:398:9  */
  assign n2053_o = n2031_o ? n2047_o : 1'b0;
  /* decoder.vhd:413:12  */
  assign n2054_o = ~clk_second_cycle_i;
  /* decoder.vhd:414:14  */
  assign n2055_o = ~int_pending_s;
  /* decoder.vhd:414:11  */
  assign n2058_o = n2055_o ? 1'b1 : 1'b0;
  /* decoder.vhd:414:11  */
  assign n2061_o = n2055_o ? 1'b0 : 1'b1;
  /* decoder.vhd:413:9  */
  assign n2063_o = n2054_o ? n2058_o : 1'b0;
  /* decoder.vhd:413:9  */
  assign n2065_o = n2054_o ? n2061_o : 1'b0;
  /* decoder.vhd:397:7  */
  assign n2067_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:422:31  */
  assign n2068_o = ~branch_taken_q;
  /* decoder.vhd:422:27  */
  assign n2069_o = n2031_o & n2068_o;
  /* decoder.vhd:423:12  */
  assign n2070_o = ~int_pending_s;
  /* decoder.vhd:422:50  */
  assign n2071_o = n2069_o & n2070_o;
  /* decoder.vhd:422:9  */
  assign n2074_o = n2071_o ? 1'b1 : 1'b0;
  /* decoder.vhd:421:7  */
  assign n2076_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:428:9  */
  assign n2079_o = n2031_o ? 1'b1 : 1'b0;
  /* decoder.vhd:427:7  */
  assign n2081_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:441:14  */
  assign n2082_o = ~clk_second_cycle_i;
  /* decoder.vhd:441:37  */
  assign n2083_o = n2082_o & assert_psen_s;
  /* decoder.vhd:442:13  */
  assign n2084_o = n2083_o | last_cycle_s;
  /* decoder.vhd:440:23  */
  assign n2085_o = ea_i & n2084_o;
  /* decoder.vhd:440:9  */
  assign n2088_o = n2085_o ? 1'b1 : 1'b0;
  /* decoder.vhd:440:9  */
  assign n2091_o = n2085_o ? 1'b1 : 1'b0;
  /* decoder.vhd:440:9  */
  assign n2094_o = n2085_o ? 1'b1 : 1'b0;
  /* decoder.vhd:439:7  */
  assign n2096_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:450:28  */
  assign n2097_o = n2031_o | last_cycle_s;
  /* decoder.vhd:449:23  */
  assign n2098_o = ea_i & n2097_o;
  /* decoder.vhd:453:12  */
  assign n2099_o = ~p2_output_exp_s;
  /* decoder.vhd:450:45  */
  assign n2100_o = n2098_o & n2099_o;
  /* decoder.vhd:455:12  */
  assign n2101_o = ~movx_first_cycle_s;
  /* decoder.vhd:453:32  */
  assign n2102_o = n2100_o & n2101_o;
  /* decoder.vhd:449:9  */
  assign n2105_o = n2102_o ? 1'b1 : 1'b0;
  /* decoder.vhd:448:7  */
  assign n2107_o = clk_mstate_i == 3'b100;
  assign n2108_o = {n2107_o, n2096_o, n2081_o, n2076_o, n2067_o};
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2110_o = 1'b0;
      5'b01000: n2110_o = 1'b0;
      5'b00100: n2110_o = 1'b0;
      5'b00010: n2110_o = 1'b0;
      5'b00001: n2110_o = n2049_o;
      default: n2110_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2113_o = 1'b0;
      5'b01000: n2113_o = n2088_o;
      5'b00100: n2113_o = 1'b0;
      5'b00010: n2113_o = 1'b0;
      5'b00001: n2113_o = 1'b0;
      default: n2113_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2116_o = 1'b0;
      5'b01000: n2116_o = n2091_o;
      5'b00100: n2116_o = 1'b0;
      5'b00010: n2116_o = 1'b0;
      5'b00001: n2116_o = 1'b0;
      default: n2116_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2119_o = n2105_o;
      5'b01000: n2119_o = n2094_o;
      5'b00100: n2119_o = 1'b0;
      5'b00010: n2119_o = 1'b0;
      5'b00001: n2119_o = n2051_o;
      default: n2119_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2122_o = 1'b0;
      5'b01000: n2122_o = 1'b0;
      5'b00100: n2122_o = 1'b0;
      5'b00010: n2122_o = 1'b0;
      5'b00001: n2122_o = n2063_o;
      default: n2122_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2125_o = 1'b0;
      5'b01000: n2125_o = 1'b0;
      5'b00100: n2125_o = 1'b0;
      5'b00010: n2125_o = 1'b0;
      5'b00001: n2125_o = n2065_o;
      default: n2125_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2128_o = 1'b0;
      5'b01000: n2128_o = 1'b0;
      5'b00100: n2128_o = 1'b0;
      5'b00010: n2128_o = n2074_o;
      5'b00001: n2128_o = 1'b0;
      default: n2128_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2131_o = 1'b0;
      5'b01000: n2131_o = 1'b0;
      5'b00100: n2131_o = n2079_o;
      5'b00010: n2131_o = 1'b0;
      5'b00001: n2131_o = 1'b0;
      default: n2131_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n2108_o)
      5'b10000: n2134_o = 1'b0;
      5'b01000: n2134_o = 1'b0;
      5'b00100: n2134_o = 1'b0;
      5'b00010: n2134_o = 1'b0;
      5'b00001: n2134_o = n2053_o;
      default: n2134_o = 1'b0;
    endcase
  /* decoder.vhd:615:5  */
  assign n2141_o = int_in_progress_s ? 1'b0 : mb_q;
  /* decoder.vhd:622:8  */
  assign n2142_o = ~clk_second_cycle_i;
  /* decoder.vhd:622:48  */
  assign n2144_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:622:31  */
  assign n2145_o = n2142_o & n2144_o;
  /* decoder.vhd:624:22  */
  assign n2146_o = opc_opcode_q[3];
  /* decoder.vhd:625:43  */
  assign n2147_o = opc_opcode_q[2:0];
  /* decoder.vhd:627:50  */
  assign n2148_o = opc_opcode_q[0];
  /* decoder.vhd:627:36  */
  assign n2150_o = {2'b00, n2148_o};
  /* decoder.vhd:624:7  */
  assign n2151_o = n2146_o ? n2147_o : n2150_o;
  assign n2153_o = n2152_o[7:3];
  /* decoder.vhd:622:5  */
  assign n2156_o = n2145_o ? 1'b1 : 1'b0;
  assign n2158_o = {n2153_o, n2151_o};
  /* decoder.vhd:622:5  */
  assign n2160_o = n2145_o ? n2158_o : 8'bX;
  /* decoder.vhd:622:5  */
  assign n2164_o = n2145_o ? 1'b1 : 1'b0;
  /* decoder.vhd:643:28  */
  assign n2166_o = opc_opcode_q[3];
  /* decoder.vhd:643:32  */
  assign n2167_o = ~n2166_o;
  /* decoder.vhd:642:44  */
  assign n2169_o = 1'b0 | n2167_o;
  /* decoder.vhd:642:13  */
  assign n2176_o = n2169_o ? 1'b1 : n2156_o;
  /* decoder.vhd:642:13  */
  assign n2179_o = n2169_o ? 1'b1 : 1'b0;
  /* decoder.vhd:642:13  */
  assign n2182_o = n2169_o ? 2'b00 : 2'b01;
  /* decoder.vhd:641:11  */
  assign n2184_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:648:11  */
  assign n2189_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:655:28  */
  assign n2193_o = opc_opcode_q[4];
  /* decoder.vhd:655:13  */
  assign n2196_o = n2193_o ? 1'b1 : 1'b0;
  /* decoder.vhd:652:11  */
  assign n2198_o = clk_mstate_i == 3'b100;
  assign n2199_o = {n2198_o, n2189_o, n2184_o};
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2202_o = 1'b1;
      3'b010: n2202_o = 1'b0;
      3'b001: n2202_o = 1'b0;
      default: n2202_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2205_o = 1'b0;
      3'b010: n2205_o = 1'b1;
      3'b001: n2205_o = 1'b0;
      default: n2205_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2208_o = 1'b1;
      3'b010: n2208_o = 1'b0;
      3'b001: n2208_o = 1'b0;
      default: n2208_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2209_o = n2156_o;
      3'b010: n2209_o = n2156_o;
      3'b001: n2209_o = n2176_o;
      default: n2209_o = n2156_o;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2212_o = 1'b0;
      3'b010: n2212_o = 1'b1;
      3'b001: n2212_o = n2179_o;
      default: n2212_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2215_o = 4'b1010;
      3'b010: n2215_o = 4'b1100;
      3'b001: n2215_o = 4'b1100;
      default: n2215_o = 4'b1100;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2217_o = n2196_o;
      3'b010: n2217_o = 1'b0;
      3'b001: n2217_o = 1'b0;
      default: n2217_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2219_o = 2'b01;
      3'b010: n2219_o = 2'b01;
      3'b001: n2219_o = n2182_o;
      default: n2219_o = 2'b01;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2221_o = alu_carry_i;
      3'b010: n2221_o = 1'b0;
      3'b001: n2221_o = 1'b0;
      default: n2221_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2224_o = 1'b1;
      3'b010: n2224_o = 1'b0;
      3'b001: n2224_o = 1'b0;
      default: n2224_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2199_o)
      3'b100: n2227_o = 1'b1;
      3'b010: n2227_o = 1'b0;
      3'b001: n2227_o = 1'b0;
      default: n2227_o = 1'b0;
    endcase
  /* decoder.vhd:638:7  */
  assign n2229_o = opc_mnemonic_s == 6'b000001;
  /* decoder.vhd:675:13  */
  assign n2231_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:682:30  */
  assign n2235_o = opc_opcode_q[4];
  /* decoder.vhd:682:15  */
  assign n2238_o = n2235_o ? 1'b1 : 1'b0;
  /* decoder.vhd:679:13  */
  assign n2240_o = clk_mstate_i == 3'b010;
  assign n2241_o = {n2240_o, n2231_o};
  /* decoder.vhd:673:11  */
  always @*
    case (n2241_o)
      2'b10: n2244_o = 1'b1;
      2'b01: n2244_o = 1'b0;
      default: n2244_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2241_o)
      2'b10: n2247_o = 1'b0;
      2'b01: n2247_o = 1'b1;
      default: n2247_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2241_o)
      2'b10: n2250_o = 1'b1;
      2'b01: n2250_o = 1'b0;
      default: n2250_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2241_o)
      2'b10: n2253_o = 4'b1010;
      2'b01: n2253_o = 4'b1100;
      default: n2253_o = 4'b1100;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2241_o)
      2'b10: n2255_o = n2238_o;
      2'b01: n2255_o = 1'b0;
      default: n2255_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2241_o)
      2'b10: n2257_o = alu_carry_i;
      2'b01: n2257_o = 1'b0;
      default: n2257_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2241_o)
      2'b10: n2260_o = 1'b1;
      2'b01: n2260_o = 1'b0;
      default: n2260_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2241_o)
      2'b10: n2263_o = 1'b1;
      2'b01: n2263_o = 1'b0;
      default: n2263_o = 1'b0;
    endcase
  /* decoder.vhd:672:9  */
  assign n2265_o = clk_second_cycle_i ? n2244_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2267_o = clk_second_cycle_i ? n2247_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2269_o = clk_second_cycle_i ? n2250_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2271_o = clk_second_cycle_i ? n2253_o : 4'b1100;
  /* decoder.vhd:672:9  */
  assign n2273_o = clk_second_cycle_i ? n2255_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2275_o = clk_second_cycle_i ? n2257_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2277_o = clk_second_cycle_i ? n2260_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2279_o = clk_second_cycle_i ? n2263_o : 1'b0;
  /* decoder.vhd:669:7  */
  assign n2281_o = opc_mnemonic_s == 6'b000010;
  /* decoder.vhd:703:28  */
  assign n2282_o = opc_opcode_q[3];
  /* decoder.vhd:703:32  */
  assign n2283_o = ~n2282_o;
  /* decoder.vhd:702:44  */
  assign n2285_o = 1'b0 | n2283_o;
  /* decoder.vhd:702:13  */
  assign n2292_o = n2285_o ? 1'b1 : n2156_o;
  /* decoder.vhd:702:13  */
  assign n2295_o = n2285_o ? 1'b1 : 1'b0;
  /* decoder.vhd:702:13  */
  assign n2298_o = n2285_o ? 2'b00 : 2'b01;
  /* decoder.vhd:701:11  */
  assign n2300_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:708:11  */
  assign n2305_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:712:11  */
  assign n2310_o = clk_mstate_i == 3'b100;
  assign n2311_o = {n2310_o, n2305_o, n2300_o};
  /* decoder.vhd:699:9  */
  always @*
    case (n2311_o)
      3'b100: n2314_o = 1'b1;
      3'b010: n2314_o = 1'b0;
      3'b001: n2314_o = 1'b0;
      default: n2314_o = 1'b0;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2311_o)
      3'b100: n2317_o = 1'b0;
      3'b010: n2317_o = 1'b1;
      3'b001: n2317_o = 1'b0;
      default: n2317_o = 1'b0;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2311_o)
      3'b100: n2320_o = 1'b1;
      3'b010: n2320_o = 1'b0;
      3'b001: n2320_o = 1'b0;
      default: n2320_o = 1'b0;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2311_o)
      3'b100: n2321_o = n2156_o;
      3'b010: n2321_o = n2156_o;
      3'b001: n2321_o = n2292_o;
      default: n2321_o = n2156_o;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2311_o)
      3'b100: n2324_o = 1'b0;
      3'b010: n2324_o = 1'b1;
      3'b001: n2324_o = n2295_o;
      default: n2324_o = 1'b0;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2311_o)
      3'b100: n2327_o = 4'b0000;
      3'b010: n2327_o = 4'b1100;
      3'b001: n2327_o = 4'b1100;
      default: n2327_o = 4'b1100;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2311_o)
      3'b100: n2329_o = 2'b01;
      3'b010: n2329_o = 2'b01;
      3'b001: n2329_o = n2298_o;
      default: n2329_o = 2'b01;
    endcase
  /* decoder.vhd:698:7  */
  assign n2331_o = opc_mnemonic_s == 6'b000011;
  /* decoder.vhd:727:13  */
  assign n2333_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:731:13  */
  assign n2338_o = clk_mstate_i == 3'b010;
  assign n2339_o = {n2338_o, n2333_o};
  /* decoder.vhd:725:11  */
  always @*
    case (n2339_o)
      2'b10: n2342_o = 1'b1;
      2'b01: n2342_o = 1'b0;
      default: n2342_o = 1'b0;
    endcase
  /* decoder.vhd:725:11  */
  always @*
    case (n2339_o)
      2'b10: n2345_o = 1'b0;
      2'b01: n2345_o = 1'b1;
      default: n2345_o = 1'b0;
    endcase
  /* decoder.vhd:725:11  */
  always @*
    case (n2339_o)
      2'b10: n2348_o = 1'b1;
      2'b01: n2348_o = 1'b0;
      default: n2348_o = 1'b0;
    endcase
  /* decoder.vhd:725:11  */
  always @*
    case (n2339_o)
      2'b10: n2351_o = 4'b0000;
      2'b01: n2351_o = 4'b1100;
      default: n2351_o = 4'b1100;
    endcase
  /* decoder.vhd:724:9  */
  assign n2353_o = clk_second_cycle_i ? n2342_o : 1'b0;
  /* decoder.vhd:724:9  */
  assign n2355_o = clk_second_cycle_i ? n2345_o : 1'b0;
  /* decoder.vhd:724:9  */
  assign n2357_o = clk_second_cycle_i ? n2348_o : 1'b0;
  /* decoder.vhd:724:9  */
  assign n2359_o = clk_second_cycle_i ? n2351_o : 4'b1100;
  /* decoder.vhd:721:7  */
  assign n2361_o = opc_mnemonic_s == 6'b000100;
  /* decoder.vhd:745:12  */
  assign n2362_o = ~clk_second_cycle_i;
  /* decoder.vhd:747:27  */
  assign n2364_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:748:28  */
  assign n2365_o = opc_opcode_q[1:0];
  /* decoder.vhd:748:41  */
  assign n2367_o = n2365_o == 2'b00;
  /* decoder.vhd:750:31  */
  assign n2368_o = opc_opcode_q[1];
  /* decoder.vhd:750:35  */
  assign n2369_o = ~n2368_o;
  /* decoder.vhd:750:13  */
  assign n2372_o = n2369_o ? 1'b1 : 1'b0;
  /* decoder.vhd:750:13  */
  assign n2375_o = n2369_o ? 1'b0 : 1'b1;
  /* decoder.vhd:750:13  */
  assign n2378_o = n2369_o ? 1'b1 : 1'b0;
  /* decoder.vhd:750:13  */
  assign n2381_o = n2369_o ? 1'b0 : 1'b1;
  /* decoder.vhd:748:13  */
  assign n2383_o = n2367_o ? 1'b0 : n2372_o;
  /* decoder.vhd:748:13  */
  assign n2385_o = n2367_o ? 1'b0 : n2375_o;
  /* decoder.vhd:748:13  */
  assign n2387_o = n2367_o ? 1'b0 : n2378_o;
  /* decoder.vhd:748:13  */
  assign n2389_o = n2367_o ? 1'b0 : n2381_o;
  /* decoder.vhd:748:13  */
  assign n2392_o = n2367_o ? 1'b1 : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2395_o = n2364_o ? 1'b1 : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2397_o = n2364_o ? n2383_o : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2399_o = n2364_o ? n2385_o : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2401_o = n2364_o ? n2387_o : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2403_o = n2364_o ? n2389_o : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2405_o = n2364_o ? n2392_o : 1'b0;
  /* decoder.vhd:765:13  */
  assign n2407_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:770:13  */
  assign n2409_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:779:30  */
  assign n2410_o = opc_opcode_q[1:0];
  /* decoder.vhd:779:43  */
  assign n2412_o = n2410_o == 2'b00;
  /* decoder.vhd:781:33  */
  assign n2413_o = opc_opcode_q[1];
  /* decoder.vhd:781:37  */
  assign n2414_o = ~n2413_o;
  /* decoder.vhd:781:15  */
  assign n2417_o = n2414_o ? 1'b1 : 1'b0;
  /* decoder.vhd:781:15  */
  assign n2420_o = n2414_o ? 1'b0 : 1'b1;
  /* decoder.vhd:779:15  */
  assign n2423_o = n2412_o ? 1'b1 : 1'b0;
  /* decoder.vhd:779:15  */
  assign n2425_o = n2412_o ? 1'b0 : n2417_o;
  /* decoder.vhd:779:15  */
  assign n2427_o = n2412_o ? 1'b0 : n2420_o;
  /* decoder.vhd:775:13  */
  assign n2429_o = clk_mstate_i == 3'b010;
  assign n2430_o = {n2429_o, n2409_o, n2407_o};
  /* decoder.vhd:762:11  */
  always @*
    case (n2430_o)
      3'b100: n2434_o = 1'b0;
      3'b010: n2434_o = 1'b1;
      3'b001: n2434_o = 1'b1;
      default: n2434_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2430_o)
      3'b100: n2438_o = 1'b1;
      3'b010: n2438_o = 1'b1;
      3'b001: n2438_o = 1'b0;
      default: n2438_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2430_o)
      3'b100: n2440_o = n2423_o;
      3'b010: n2440_o = 1'b0;
      3'b001: n2440_o = 1'b0;
      default: n2440_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2430_o)
      3'b100: n2442_o = n2425_o;
      3'b010: n2442_o = 1'b0;
      3'b001: n2442_o = 1'b0;
      default: n2442_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2430_o)
      3'b100: n2444_o = n2427_o;
      3'b010: n2444_o = 1'b0;
      3'b001: n2444_o = 1'b0;
      default: n2444_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2430_o)
      3'b100: n2447_o = 4'b0000;
      3'b010: n2447_o = 4'b1100;
      3'b001: n2447_o = 4'b1100;
      default: n2447_o = 4'b1100;
    endcase
  /* decoder.vhd:745:9  */
  assign n2449_o = n2362_o ? 1'b0 : n2434_o;
  /* decoder.vhd:745:9  */
  assign n2451_o = n2362_o ? n2395_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2453_o = n2362_o ? 1'b0 : n2438_o;
  /* decoder.vhd:745:9  */
  assign n2455_o = n2362_o ? 1'b0 : n2440_o;
  /* decoder.vhd:745:9  */
  assign n2457_o = n2362_o ? 1'b0 : n2442_o;
  /* decoder.vhd:745:9  */
  assign n2459_o = n2362_o ? n2397_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2461_o = n2362_o ? 1'b0 : n2444_o;
  /* decoder.vhd:745:9  */
  assign n2463_o = n2362_o ? n2399_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2465_o = n2362_o ? 4'b1100 : n2447_o;
  /* decoder.vhd:745:9  */
  assign n2467_o = n2362_o ? n2401_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2469_o = n2362_o ? n2403_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2471_o = n2362_o ? n2405_o : 1'b0;
  /* decoder.vhd:742:7  */
  assign n2473_o = opc_mnemonic_s == 6'b000101;
  /* decoder.vhd:798:12  */
  assign n2474_o = ~clk_second_cycle_i;
  /* decoder.vhd:811:18  */
  assign n2475_o = ~int_pending_s;
  /* decoder.vhd:811:15  */
  assign n2478_o = n2475_o ? 1'b1 : 1'b0;
  /* decoder.vhd:802:13  */
  assign n2480_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:816:13  */
  assign n2482_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:822:13  */
  assign n2484_o = clk_mstate_i == 3'b100;
  assign n2485_o = {n2484_o, n2482_o, n2480_o};
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2488_o = 1'b1;
      3'b010: n2488_o = n2156_o;
      3'b001: n2488_o = 1'b1;
      default: n2488_o = n2156_o;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2491_o = 1'b0;
      3'b010: n2491_o = 1'b1;
      3'b001: n2491_o = 1'b0;
      default: n2491_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2494_o = 1'b1;
      3'b010: n2494_o = 1'b0;
      3'b001: n2494_o = 1'b0;
      default: n2494_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2497_o = 1'b1;
      3'b010: n2497_o = 1'b0;
      3'b001: n2497_o = 1'b0;
      default: n2497_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2500_o = 1'b0;
      3'b010: n2500_o = 1'b0;
      3'b001: n2500_o = 1'b1;
      default: n2500_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2504_o = 2'b11;
      3'b010: n2504_o = 2'b01;
      3'b001: n2504_o = 2'b10;
      default: n2504_o = 2'b01;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2507_o = 1'b1;
      3'b010: n2507_o = 1'b0;
      3'b001: n2507_o = 1'b0;
      default: n2507_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2509_o = 1'b0;
      3'b010: n2509_o = 1'b0;
      3'b001: n2509_o = n2478_o;
      default: n2509_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2485_o)
      3'b100: n2513_o = 1'b1;
      3'b010: n2513_o = 1'b1;
      3'b001: n2513_o = 1'b0;
      default: n2513_o = 1'b0;
    endcase
  /* decoder.vhd:845:17  */
  assign n2520_o = tim_int_s ? 1'b0 : 1'b1;
  assign n2521_o = n2515_o[2];
  /* decoder.vhd:845:17  */
  assign n2522_o = tim_int_s ? 1'b1 : n2521_o;
  assign n2523_o = n2515_o[7:3];
  /* decoder.vhd:841:15  */
  assign n2525_o = int_pending_s ? n2520_o : 1'b0;
  assign n2526_o = {n2523_o, n2522_o, 2'b11};
  /* decoder.vhd:841:15  */
  assign n2527_o = int_pending_s ? n2526_o : n2160_o;
  /* decoder.vhd:841:15  */
  assign n2529_o = int_pending_s ? 1'b1 : n2164_o;
  /* decoder.vhd:838:13  */
  assign n2531_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:856:18  */
  assign n2532_o = ~int_pending_s;
  /* decoder.vhd:858:46  */
  assign n2534_o = {4'b0000, n2141_o};
  /* decoder.vhd:858:67  */
  assign n2535_o = opc_opcode_q[7:5];
  /* decoder.vhd:858:53  */
  assign n2536_o = {n2534_o, n2535_o};
  /* decoder.vhd:856:15  */
  assign n2538_o = n2532_o ? n2536_o : 8'b00000000;
  /* decoder.vhd:856:15  */
  assign n2541_o = n2532_o ? 1'b0 : 1'b1;
  /* decoder.vhd:853:13  */
  assign n2543_o = clk_mstate_i == 3'b001;
  assign n2544_o = {n2543_o, n2531_o};
  /* decoder.vhd:836:11  */
  always @*
    case (n2544_o)
      2'b10: n2546_o = 1'b0;
      2'b01: n2546_o = n2525_o;
      default: n2546_o = 1'b0;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2544_o)
      2'b10: n2549_o = 1'b0;
      2'b01: n2549_o = 1'b1;
      default: n2549_o = 1'b0;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2544_o)
      2'b10: n2552_o = 1'b1;
      2'b01: n2552_o = 1'b0;
      default: n2552_o = 1'b0;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2544_o)
      2'b10: n2555_o = 1'b0;
      2'b01: n2555_o = 1'b1;
      default: n2555_o = 1'b0;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2544_o)
      2'b10: n2556_o = n2538_o;
      2'b01: n2556_o = n2527_o;
      default: n2556_o = n2160_o;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2544_o)
      2'b10: n2558_o = 1'b1;
      2'b01: n2558_o = n2529_o;
      default: n2558_o = n2164_o;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2544_o)
      2'b10: n2560_o = n2541_o;
      2'b01: n2560_o = 1'b0;
      default: n2560_o = 1'b0;
    endcase
  /* decoder.vhd:798:9  */
  assign n2562_o = n2474_o ? 1'b0 : n2546_o;
  /* decoder.vhd:798:9  */
  assign n2563_o = n2474_o ? n2488_o : n2156_o;
  /* decoder.vhd:798:9  */
  assign n2565_o = n2474_o ? 1'b0 : n2549_o;
  /* decoder.vhd:798:9  */
  assign n2567_o = n2474_o ? n2491_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2569_o = n2474_o ? 1'b0 : n2552_o;
  /* decoder.vhd:798:9  */
  assign n2571_o = n2474_o ? n2494_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2573_o = n2474_o ? n2497_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2575_o = n2474_o ? n2500_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2577_o = n2474_o ? n2504_o : 2'b01;
  /* decoder.vhd:798:9  */
  assign n2579_o = n2474_o ? n2507_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2581_o = n2474_o ? 1'b0 : n2555_o;
  /* decoder.vhd:798:9  */
  assign n2583_o = n2474_o ? n2509_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2584_o = n2474_o ? n2160_o : n2556_o;
  /* decoder.vhd:798:9  */
  assign n2585_o = n2474_o ? n2164_o : n2558_o;
  /* decoder.vhd:798:9  */
  assign n2587_o = n2474_o ? n2513_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2589_o = n2474_o ? 1'b0 : n2560_o;
  /* decoder.vhd:795:7  */
  assign n2591_o = opc_mnemonic_s == 6'b000110;
  /* decoder.vhd:875:25  */
  assign n2593_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:875:9  */
  assign n2596_o = n2593_o ? 1'b1 : 1'b0;
  /* decoder.vhd:875:9  */
  assign n2599_o = n2593_o ? 1'b1 : 1'b0;
  /* decoder.vhd:875:9  */
  assign n2602_o = n2593_o ? 4'b0100 : 4'b1100;
  /* decoder.vhd:873:7  */
  assign n2604_o = opc_mnemonic_s == 6'b000111;
  /* decoder.vhd:884:25  */
  assign n2606_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:884:9  */
  assign n2609_o = n2606_o ? 1'b1 : 1'b0;
  /* decoder.vhd:882:7  */
  assign n2611_o = opc_mnemonic_s == 6'b001000;
  /* decoder.vhd:892:25  */
  assign n2613_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:893:26  */
  assign n2614_o = opc_opcode_q[5];
  /* decoder.vhd:893:30  */
  assign n2615_o = ~n2614_o;
  /* decoder.vhd:893:11  */
  assign n2618_o = n2615_o ? 1'b1 : 1'b0;
  /* decoder.vhd:893:11  */
  assign n2621_o = n2615_o ? 1'b0 : 1'b1;
  /* decoder.vhd:892:9  */
  assign n2623_o = n2613_o ? n2618_o : 1'b0;
  /* decoder.vhd:892:9  */
  assign n2625_o = n2613_o ? n2621_o : 1'b0;
  /* decoder.vhd:890:7  */
  assign n2627_o = opc_mnemonic_s == 6'b001001;
  /* decoder.vhd:905:25  */
  assign n2629_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:905:9  */
  assign n2632_o = n2629_o ? 1'b1 : 1'b0;
  /* decoder.vhd:905:9  */
  assign n2635_o = n2629_o ? 1'b1 : 1'b0;
  /* decoder.vhd:905:9  */
  assign n2638_o = n2629_o ? 4'b0011 : 4'b1100;
  /* decoder.vhd:903:7  */
  assign n2640_o = opc_mnemonic_s == 6'b001010;
  /* decoder.vhd:914:25  */
  assign n2642_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:915:33  */
  assign n2643_o = ~psw_carry_i;
  /* decoder.vhd:914:9  */
  assign n2645_o = n2642_o ? n2643_o : 1'b0;
  /* decoder.vhd:914:9  */
  assign n2648_o = n2642_o ? 1'b1 : 1'b0;
  /* decoder.vhd:912:7  */
  assign n2650_o = opc_mnemonic_s == 6'b001011;
  /* decoder.vhd:922:25  */
  assign n2652_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:923:26  */
  assign n2653_o = opc_opcode_q[5];
  /* decoder.vhd:923:30  */
  assign n2654_o = ~n2653_o;
  /* decoder.vhd:924:35  */
  assign n2655_o = ~psw_f0_i;
  /* decoder.vhd:923:11  */
  assign n2657_o = n2654_o ? n2655_o : 1'b0;
  /* decoder.vhd:923:11  */
  assign n2660_o = n2654_o ? 1'b1 : 1'b0;
  /* decoder.vhd:923:11  */
  assign n2663_o = n2654_o ? 1'b0 : 1'b1;
  /* decoder.vhd:922:9  */
  assign n2665_o = n2652_o ? n2657_o : 1'b0;
  /* decoder.vhd:922:9  */
  assign n2667_o = n2652_o ? n2660_o : 1'b0;
  /* decoder.vhd:922:9  */
  assign n2669_o = n2652_o ? n2663_o : 1'b0;
  /* decoder.vhd:920:7  */
  assign n2671_o = opc_mnemonic_s == 6'b001100;
  /* decoder.vhd:938:11  */
  assign n2673_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:944:38  */
  assign n2674_o = psw_aux_carry_i | alu_da_overflow_i;
  /* decoder.vhd:944:13  */
  assign n2677_o = n2674_o ? 1'b1 : 1'b0;
  /* decoder.vhd:944:13  */
  assign n2680_o = n2674_o ? 1'b1 : 1'b0;
  /* decoder.vhd:943:11  */
  assign n2682_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:958:13  */
  assign n2685_o = alu_da_overflow_i ? 4'b1010 : 4'b1100;
  /* decoder.vhd:958:13  */
  assign n2687_o = alu_da_overflow_i ? alu_carry_i : 1'b0;
  /* decoder.vhd:955:11  */
  assign n2689_o = clk_mstate_i == 3'b100;
  assign n2690_o = {n2689_o, n2682_o, n2673_o};
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2693_o = 1'b1;
      3'b010: n2693_o = 1'b0;
      3'b001: n2693_o = 1'b0;
      default: n2693_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2695_o = 1'b0;
      3'b010: n2695_o = n2677_o;
      3'b001: n2695_o = 1'b0;
      default: n2695_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2698_o = 1'b1;
      3'b010: n2698_o = n2680_o;
      3'b001: n2698_o = 1'b0;
      default: n2698_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2700_o = n2685_o;
      3'b010: n2700_o = 4'b1010;
      3'b001: n2700_o = 4'b1010;
      default: n2700_o = 4'b1010;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2704_o = 1'b1;
      3'b010: n2704_o = 1'b0;
      3'b001: n2704_o = 1'b0;
      default: n2704_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2707_o = 1'b0;
      3'b010: n2707_o = 1'b0;
      3'b001: n2707_o = 1'b1;
      default: n2707_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2710_o = 1'b0;
      3'b010: n2710_o = 1'b1;
      3'b001: n2710_o = 1'b0;
      default: n2710_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2712_o = n2687_o;
      3'b010: n2712_o = 1'b0;
      3'b001: n2712_o = 1'b0;
      default: n2712_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2690_o)
      3'b100: n2715_o = 1'b1;
      3'b010: n2715_o = 1'b0;
      3'b001: n2715_o = 1'b0;
      default: n2715_o = 1'b0;
    endcase
  /* decoder.vhd:933:7  */
  assign n2717_o = opc_mnemonic_s == 6'b001101;
  /* decoder.vhd:978:28  */
  assign n2718_o = opc_opcode_q[6];
  /* decoder.vhd:978:13  */
  assign n2721_o = n2718_o ? 1'b1 : 1'b0;
  /* decoder.vhd:978:13  */
  assign n2724_o = n2718_o ? 1'b1 : 1'b0;
  /* decoder.vhd:976:11  */
  assign n2726_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:987:28  */
  assign n2727_o = opc_opcode_q[6];
  /* decoder.vhd:987:32  */
  assign n2728_o = ~n2727_o;
  /* decoder.vhd:987:13  */
  assign n2731_o = n2728_o ? 1'b1 : 1'b0;
  /* decoder.vhd:987:13  */
  assign n2734_o = n2728_o ? 1'b0 : 1'b1;
  /* decoder.vhd:983:11  */
  assign n2736_o = clk_mstate_i == 3'b100;
  assign n2737_o = {n2736_o, n2726_o};
  /* decoder.vhd:975:9  */
  always @*
    case (n2737_o)
      2'b10: n2739_o = n2731_o;
      2'b01: n2739_o = 1'b0;
      default: n2739_o = 1'b0;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2737_o)
      2'b10: n2741_o = 1'b0;
      2'b01: n2741_o = n2721_o;
      default: n2741_o = 1'b0;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2737_o)
      2'b10: n2744_o = 1'b1;
      2'b01: n2744_o = 1'b0;
      default: n2744_o = 1'b0;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2737_o)
      2'b10: n2746_o = 1'b0;
      2'b01: n2746_o = n2724_o;
      default: n2746_o = 1'b0;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2737_o)
      2'b10: n2749_o = 4'b1000;
      2'b01: n2749_o = 4'b1100;
      default: n2749_o = 4'b1100;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2737_o)
      2'b10: n2751_o = n2734_o;
      2'b01: n2751_o = 1'b0;
      default: n2751_o = 1'b0;
    endcase
  /* decoder.vhd:974:7  */
  assign n2753_o = opc_mnemonic_s == 6'b001110;
  /* decoder.vhd:1002:25  */
  assign n2755_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1003:26  */
  assign n2756_o = opc_opcode_q[4];
  /* decoder.vhd:1003:11  */
  assign n2759_o = n2756_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1003:11  */
  assign n2762_o = n2756_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1002:9  */
  assign n2764_o = n2755_o ? n2759_o : 1'b0;
  /* decoder.vhd:1002:9  */
  assign n2766_o = n2755_o ? n2762_o : 1'b0;
  /* decoder.vhd:1001:7  */
  assign n2768_o = opc_mnemonic_s == 6'b001111;
  /* decoder.vhd:1012:25  */
  assign n2770_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1013:26  */
  assign n2771_o = opc_opcode_q[4];
  /* decoder.vhd:1013:11  */
  assign n2774_o = n2771_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1013:11  */
  assign n2777_o = n2771_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1012:9  */
  assign n2779_o = n2770_o ? n2774_o : 1'b0;
  /* decoder.vhd:1012:9  */
  assign n2781_o = n2770_o ? n2777_o : 1'b0;
  /* decoder.vhd:1011:7  */
  assign n2783_o = opc_mnemonic_s == 6'b010000;
  /* decoder.vhd:1024:12  */
  assign n2784_o = ~clk_second_cycle_i;
  /* decoder.vhd:1027:13  */
  assign n2786_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1033:13  */
  assign n2789_o = clk_mstate_i == 3'b100;
  assign n2790_o = {n2789_o, n2786_o};
  /* decoder.vhd:1025:11  */
  always @*
    case (n2790_o)
      2'b10: n2793_o = 1'b0;
      2'b01: n2793_o = 1'b1;
      default: n2793_o = 1'b0;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2790_o)
      2'b10: n2796_o = 1'b1;
      2'b01: n2796_o = 1'b0;
      default: n2796_o = 1'b0;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2790_o)
      2'b10: n2799_o = 1'b0;
      2'b01: n2799_o = 1'b1;
      default: n2799_o = 1'b0;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2790_o)
      2'b10: n2802_o = 4'b1000;
      2'b01: n2802_o = 4'b1100;
      default: n2802_o = 4'b1100;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2790_o)
      2'b10: n2805_o = 1'b1;
      2'b01: n2805_o = 1'b0;
      default: n2805_o = 1'b0;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2790_o)
      2'b10: n2808_o = 4'b0001;
      2'b01: n2808_o = 4'b0000;
      default: n2808_o = 4'b0000;
    endcase
  assign n2809_o = opc_opcode_q[5];
  /* decoder.vhd:1025:11  */
  always @*
    case (n2790_o)
      2'b10: n2810_o = 1'b0;
      2'b01: n2810_o = n2809_o;
      default: n2810_o = n2809_o;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2790_o)
      2'b10: n2813_o = 1'b1;
      2'b01: n2813_o = 1'b0;
      default: n2813_o = 1'b0;
    endcase
  /* decoder.vhd:1050:27  */
  assign n2815_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1050:37  */
  assign n2816_o = n2815_o & cnd_take_branch_i;
  /* decoder.vhd:1050:11  */
  assign n2822_o = n2816_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1050:11  */
  assign n2825_o = n2816_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2827_o = n2784_o ? n2793_o : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2829_o = n2784_o ? n2796_o : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2831_o = n2784_o ? n2799_o : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2833_o = n2784_o ? 1'b0 : n2822_o;
  /* decoder.vhd:1024:9  */
  assign n2835_o = n2784_o ? n2802_o : 4'b1100;
  /* decoder.vhd:1024:9  */
  assign n2837_o = n2784_o ? n2805_o : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2839_o = n2784_o ? n2808_o : 4'b0000;
  assign n2840_o = opc_opcode_q[5];
  /* decoder.vhd:1024:9  */
  assign n2841_o = n2784_o ? n2810_o : n2840_o;
  /* decoder.vhd:1024:9  */
  assign n2843_o = n2784_o ? 1'b0 : n2825_o;
  /* decoder.vhd:1024:9  */
  assign n2845_o = n2784_o ? n2813_o : 1'b0;
  /* decoder.vhd:1021:7  */
  assign n2847_o = opc_mnemonic_s == 6'b010001;
  /* decoder.vhd:1058:25  */
  assign n2849_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1059:26  */
  assign n2850_o = opc_opcode_q[4];
  /* decoder.vhd:1059:30  */
  assign n2851_o = ~n2850_o;
  /* decoder.vhd:1059:11  */
  assign n2854_o = n2851_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1059:11  */
  assign n2857_o = n2851_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1058:9  */
  assign n2859_o = n2849_o ? n2854_o : 1'b0;
  /* decoder.vhd:1058:9  */
  assign n2861_o = n2849_o ? n2857_o : 1'b0;
  /* decoder.vhd:1057:7  */
  assign n2863_o = opc_mnemonic_s == 6'b111110;
  /* decoder.vhd:1068:25  */
  assign n2865_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1068:9  */
  assign n2868_o = n2865_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1067:7  */
  assign n2870_o = opc_mnemonic_s == 6'b010010;
  /* decoder.vhd:1075:48  */
  assign n2872_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1075:31  */
  assign n2873_o = clk_second_cycle_i & n2872_o;
  /* decoder.vhd:1078:26  */
  assign n2874_o = opc_opcode_q[1];
  /* decoder.vhd:1078:30  */
  assign n2875_o = ~n2874_o;
  /* decoder.vhd:1078:11  */
  assign n2878_o = n2875_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1078:11  */
  assign n2881_o = n2875_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1075:9  */
  assign n2884_o = n2873_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1075:9  */
  assign n2886_o = n2873_o ? n2878_o : 1'b0;
  /* decoder.vhd:1075:9  */
  assign n2888_o = n2873_o ? n2881_o : 1'b0;
  /* decoder.vhd:1073:7  */
  assign n2890_o = opc_mnemonic_s == 6'b010011;
  /* decoder.vhd:1088:25  */
  assign n2892_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1088:9  */
  assign n2895_o = n2892_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1088:9  */
  assign n2898_o = n2892_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1086:7  */
  assign n2900_o = opc_mnemonic_s == 6'b111010;
  /* decoder.vhd:1099:48  */
  assign n2902_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1099:31  */
  assign n2903_o = clk_second_cycle_i & n2902_o;
  /* decoder.vhd:1099:9  */
  assign n2906_o = n2903_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1099:9  */
  assign n2909_o = n2903_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1095:7  */
  assign n2911_o = opc_mnemonic_s == 6'b010101;
  /* decoder.vhd:1111:28  */
  assign n2912_o = opc_opcode_q[3];
  /* decoder.vhd:1111:32  */
  assign n2913_o = ~n2912_o;
  /* decoder.vhd:1110:44  */
  assign n2915_o = 1'b0 | n2913_o;
  /* decoder.vhd:1110:13  */
  assign n2922_o = n2915_o ? 1'b1 : n2156_o;
  /* decoder.vhd:1110:13  */
  assign n2925_o = n2915_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1110:13  */
  assign n2928_o = n2915_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1109:11  */
  assign n2930_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1117:28  */
  assign n2931_o = opc_opcode_q[3:2];
  /* decoder.vhd:1117:41  */
  assign n2933_o = n2931_o != 2'b01;
  /* decoder.vhd:1117:13  */
  assign n2936_o = n2933_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1117:13  */
  assign n2939_o = n2933_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1115:11  */
  assign n2941_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1126:28  */
  assign n2942_o = opc_opcode_q[3:2];
  /* decoder.vhd:1126:41  */
  assign n2944_o = n2942_o == 2'b01;
  /* decoder.vhd:1126:13  */
  assign n2947_o = n2944_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1126:13  */
  assign n2950_o = n2944_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1122:11  */
  assign n2952_o = clk_mstate_i == 3'b100;
  assign n2953_o = {n2952_o, n2941_o, n2930_o};
  /* decoder.vhd:1107:9  */
  always @*
    case (n2953_o)
      3'b100: n2955_o = n2947_o;
      3'b010: n2955_o = 1'b0;
      3'b001: n2955_o = 1'b0;
      default: n2955_o = 1'b0;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2953_o)
      3'b100: n2957_o = 1'b0;
      3'b010: n2957_o = n2936_o;
      3'b001: n2957_o = 1'b0;
      default: n2957_o = 1'b0;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2953_o)
      3'b100: n2960_o = 1'b1;
      3'b010: n2960_o = 1'b0;
      3'b001: n2960_o = 1'b0;
      default: n2960_o = 1'b0;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2953_o)
      3'b100: n2961_o = n2156_o;
      3'b010: n2961_o = n2156_o;
      3'b001: n2961_o = n2922_o;
      default: n2961_o = n2156_o;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2953_o)
      3'b100: n2963_o = 1'b0;
      3'b010: n2963_o = n2939_o;
      3'b001: n2963_o = n2925_o;
      default: n2963_o = 1'b0;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2953_o)
      3'b100: n2966_o = 4'b1001;
      3'b010: n2966_o = 4'b1100;
      3'b001: n2966_o = 4'b1100;
      default: n2966_o = 4'b1100;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2953_o)
      3'b100: n2968_o = 2'b01;
      3'b010: n2968_o = 2'b01;
      3'b001: n2968_o = n2928_o;
      default: n2968_o = 2'b01;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2953_o)
      3'b100: n2970_o = n2950_o;
      3'b010: n2970_o = 1'b0;
      3'b001: n2970_o = 1'b0;
      default: n2970_o = 1'b0;
    endcase
  /* decoder.vhd:1106:7  */
  assign n2972_o = opc_mnemonic_s == 6'b010100;
  /* decoder.vhd:1144:12  */
  assign n2973_o = ~clk_second_cycle_i;
  /* decoder.vhd:1146:27  */
  assign n2975_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1146:11  */
  assign n2978_o = n2975_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1146:11  */
  assign n2981_o = n2975_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1155:27  */
  assign n2983_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1155:37  */
  assign n2984_o = n2983_o & cnd_take_branch_i;
  /* decoder.vhd:1155:11  */
  assign n2990_o = n2984_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1155:11  */
  assign n2993_o = n2984_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1144:9  */
  assign n2995_o = n2973_o ? n2978_o : 1'b0;
  /* decoder.vhd:1144:9  */
  assign n2997_o = n2973_o ? 1'b0 : n2990_o;
  /* decoder.vhd:1144:9  */
  assign n2999_o = n2973_o ? n2981_o : 1'b0;
  /* decoder.vhd:1144:9  */
  assign n3001_o = n2973_o ? 1'b0 : n2993_o;
  /* decoder.vhd:1140:7  */
  assign n3003_o = opc_mnemonic_s == 6'b010110;
  /* decoder.vhd:1166:12  */
  assign n3004_o = ~clk_second_cycle_i;
  /* decoder.vhd:1168:27  */
  assign n3006_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1170:48  */
  assign n3007_o = opc_opcode_q[4];
  /* decoder.vhd:1168:11  */
  assign n3010_o = n3006_o ? 1'b1 : 1'b0;
  assign n3011_o = opc_opcode_q[5];
  /* decoder.vhd:1166:9  */
  assign n3012_o = n3030_o ? n3007_o : n3011_o;
  /* decoder.vhd:1176:27  */
  assign n3014_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1176:37  */
  assign n3015_o = n3014_o & cnd_take_branch_i;
  /* decoder.vhd:1176:11  */
  assign n3021_o = n3015_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1176:11  */
  assign n3024_o = n3015_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1166:9  */
  assign n3026_o = n3004_o ? 1'b0 : n3021_o;
  /* decoder.vhd:1166:9  */
  assign n3028_o = n3004_o ? n3010_o : 1'b0;
  /* decoder.vhd:1166:9  */
  assign n3030_o = n3004_o & n3006_o;
  /* decoder.vhd:1166:9  */
  assign n3032_o = n3004_o ? 1'b0 : n3024_o;
  /* decoder.vhd:1162:7  */
  assign n3034_o = opc_mnemonic_s == 6'b010111;
  /* decoder.vhd:1186:12  */
  assign n3035_o = ~clk_second_cycle_i;
  /* decoder.vhd:1188:27  */
  assign n3037_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1190:28  */
  assign n3038_o = opc_opcode_q[7];
  /* decoder.vhd:1190:13  */
  assign n3041_o = n3038_o ? 4'b0011 : 4'b0100;
  /* decoder.vhd:1188:11  */
  assign n3044_o = n3037_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1188:11  */
  assign n3046_o = n3037_o ? n3041_o : 4'b0000;
  /* decoder.vhd:1203:27  */
  assign n3048_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1203:37  */
  assign n3049_o = n3048_o & cnd_take_branch_i;
  /* decoder.vhd:1203:11  */
  assign n3055_o = n3049_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1203:11  */
  assign n3058_o = n3049_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1186:9  */
  assign n3060_o = n3035_o ? 1'b0 : n3055_o;
  /* decoder.vhd:1186:9  */
  assign n3062_o = n3035_o ? n3044_o : 1'b0;
  /* decoder.vhd:1186:9  */
  assign n3064_o = n3035_o ? n3046_o : 4'b0000;
  /* decoder.vhd:1186:9  */
  assign n3066_o = n3035_o ? 1'b0 : n3058_o;
  /* decoder.vhd:1183:7  */
  assign n3068_o = opc_mnemonic_s == 6'b011000;
  /* decoder.vhd:1217:13  */
  assign n3070_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1223:40  */
  assign n3072_o = {4'b0000, n2141_o};
  /* decoder.vhd:1223:61  */
  assign n3073_o = opc_opcode_q[7:5];
  /* decoder.vhd:1223:47  */
  assign n3074_o = {n3072_o, n3073_o};
  /* decoder.vhd:1222:13  */
  assign n3076_o = clk_mstate_i == 3'b001;
  assign n3077_o = {n3076_o, n3070_o};
  /* decoder.vhd:1215:11  */
  always @*
    case (n3077_o)
      2'b10: n3080_o = 1'b0;
      2'b01: n3080_o = 1'b1;
      default: n3080_o = 1'b0;
    endcase
  /* decoder.vhd:1215:11  */
  always @*
    case (n3077_o)
      2'b10: n3083_o = 1'b1;
      2'b01: n3083_o = 1'b0;
      default: n3083_o = 1'b0;
    endcase
  /* decoder.vhd:1215:11  */
  always @*
    case (n3077_o)
      2'b10: n3086_o = 1'b0;
      2'b01: n3086_o = 1'b1;
      default: n3086_o = 1'b0;
    endcase
  /* decoder.vhd:1215:11  */
  always @*
    case (n3077_o)
      2'b10: n3087_o = n3074_o;
      2'b01: n3087_o = n2160_o;
      default: n3087_o = n2160_o;
    endcase
  /* decoder.vhd:1215:11  */
  always @*
    case (n3077_o)
      2'b10: n3089_o = 1'b1;
      2'b01: n3089_o = n2164_o;
      default: n3089_o = n2164_o;
    endcase
  /* decoder.vhd:1214:9  */
  assign n3091_o = clk_second_cycle_i ? n3080_o : 1'b0;
  /* decoder.vhd:1214:9  */
  assign n3093_o = clk_second_cycle_i ? n3083_o : 1'b0;
  /* decoder.vhd:1214:9  */
  assign n3095_o = clk_second_cycle_i ? n3086_o : 1'b0;
  /* decoder.vhd:1214:9  */
  assign n3096_o = clk_second_cycle_i ? n3087_o : n2160_o;
  /* decoder.vhd:1214:9  */
  assign n3097_o = clk_second_cycle_i ? n3089_o : n2164_o;
  /* decoder.vhd:1211:7  */
  assign n3099_o = opc_mnemonic_s == 6'b011001;
  /* decoder.vhd:1238:12  */
  assign n3100_o = ~clk_second_cycle_i;
  /* decoder.vhd:1241:27  */
  assign n3102_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1241:11  */
  assign n3105_o = n3102_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1241:11  */
  assign n3108_o = n3102_o ? 2'b01 : 2'b00;
  /* decoder.vhd:1247:27  */
  assign n3110_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1247:11  */
  assign n3113_o = n3110_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1247:11  */
  assign n3116_o = n3110_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1238:9  */
  assign n3118_o = n3100_o ? n3105_o : 1'b0;
  /* decoder.vhd:1238:9  */
  assign n3120_o = n3100_o ? 1'b0 : n3113_o;
  /* decoder.vhd:1238:9  */
  assign n3122_o = n3100_o ? n3108_o : 2'b00;
  /* decoder.vhd:1238:9  */
  assign n3124_o = n3100_o ? 1'b0 : n3116_o;
  /* decoder.vhd:1235:7  */
  assign n3126_o = opc_mnemonic_s == 6'b011010;
  /* decoder.vhd:1260:12  */
  assign n3127_o = ~clk_second_cycle_i;
  /* decoder.vhd:1262:27  */
  assign n3129_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1262:11  */
  assign n3132_o = n3129_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1269:27  */
  assign n3134_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1269:37  */
  assign n3135_o = n3134_o & cnd_take_branch_i;
  /* decoder.vhd:1269:11  */
  assign n3141_o = n3135_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1269:11  */
  assign n3144_o = n3135_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1260:9  */
  assign n3146_o = n3127_o ? 1'b0 : n3141_o;
  /* decoder.vhd:1260:9  */
  assign n3148_o = n3127_o ? n3132_o : 1'b0;
  /* decoder.vhd:1260:9  */
  assign n3150_o = n3127_o ? 1'b0 : n3144_o;
  /* decoder.vhd:1256:7  */
  assign n3152_o = opc_mnemonic_s == 6'b011011;
  /* decoder.vhd:1280:12  */
  assign n3153_o = ~clk_second_cycle_i;
  /* decoder.vhd:1282:27  */
  assign n3155_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1282:11  */
  assign n3158_o = n3155_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1289:27  */
  assign n3160_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1289:37  */
  assign n3161_o = n3160_o & cnd_take_branch_i;
  /* decoder.vhd:1289:11  */
  assign n3167_o = n3161_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1289:11  */
  assign n3170_o = n3161_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1280:9  */
  assign n3172_o = n3153_o ? 1'b0 : n3167_o;
  /* decoder.vhd:1280:9  */
  assign n3174_o = n3153_o ? n3158_o : 1'b0;
  /* decoder.vhd:1280:9  */
  assign n3176_o = n3153_o ? 1'b0 : n3170_o;
  /* decoder.vhd:1276:7  */
  assign n3178_o = opc_mnemonic_s == 6'b111100;
  /* decoder.vhd:1300:12  */
  assign n3179_o = ~clk_second_cycle_i;
  /* decoder.vhd:1302:27  */
  assign n3181_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1302:11  */
  assign n3184_o = n3181_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1309:27  */
  assign n3186_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1309:37  */
  assign n3187_o = n3186_o & cnd_take_branch_i;
  /* decoder.vhd:1309:11  */
  assign n3193_o = n3187_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1309:11  */
  assign n3196_o = n3187_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1300:9  */
  assign n3198_o = n3179_o ? 1'b0 : n3193_o;
  /* decoder.vhd:1300:9  */
  assign n3200_o = n3179_o ? n3184_o : 1'b0;
  /* decoder.vhd:1300:9  */
  assign n3202_o = n3179_o ? 1'b0 : n3196_o;
  /* decoder.vhd:1296:7  */
  assign n3204_o = opc_mnemonic_s == 6'b111101;
  /* decoder.vhd:1318:24  */
  assign n3205_o = opc_opcode_q[6];
  /* decoder.vhd:1318:28  */
  assign n3206_o = ~n3205_o;
  /* decoder.vhd:1318:9  */
  assign n3209_o = n3206_o ? 4'b0110 : 4'b0111;
  /* decoder.vhd:1324:12  */
  assign n3210_o = ~clk_second_cycle_i;
  /* decoder.vhd:1326:27  */
  assign n3212_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1328:48  */
  assign n3213_o = opc_opcode_q[4];
  /* decoder.vhd:1326:11  */
  assign n3216_o = n3212_o ? 1'b1 : 1'b0;
  assign n3217_o = opc_opcode_q[5];
  /* decoder.vhd:1324:9  */
  assign n3218_o = n3236_o ? n3213_o : n3217_o;
  /* decoder.vhd:1334:27  */
  assign n3220_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1334:37  */
  assign n3221_o = n3220_o & cnd_take_branch_i;
  /* decoder.vhd:1334:11  */
  assign n3227_o = n3221_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1334:11  */
  assign n3230_o = n3221_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1324:9  */
  assign n3232_o = n3210_o ? 1'b0 : n3227_o;
  /* decoder.vhd:1324:9  */
  assign n3234_o = n3210_o ? n3216_o : 1'b0;
  /* decoder.vhd:1324:9  */
  assign n3236_o = n3210_o & n3212_o;
  /* decoder.vhd:1324:9  */
  assign n3238_o = n3210_o ? 1'b0 : n3230_o;
  /* decoder.vhd:1316:7  */
  assign n3240_o = opc_mnemonic_s == 6'b011100;
  /* decoder.vhd:1345:12  */
  assign n3241_o = ~clk_second_cycle_i;
  /* decoder.vhd:1347:27  */
  assign n3243_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1347:11  */
  assign n3246_o = n3243_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1347:11  */
  assign n3249_o = n3243_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1355:27  */
  assign n3251_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1355:37  */
  assign n3252_o = n3251_o & cnd_take_branch_i;
  /* decoder.vhd:1355:11  */
  assign n3258_o = n3252_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1355:11  */
  assign n3261_o = n3252_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1345:9  */
  assign n3263_o = n3241_o ? 1'b0 : n3258_o;
  /* decoder.vhd:1345:9  */
  assign n3265_o = n3241_o ? n3246_o : 1'b0;
  /* decoder.vhd:1345:9  */
  assign n3267_o = n3241_o ? 1'b0 : n3261_o;
  /* decoder.vhd:1345:9  */
  assign n3269_o = n3241_o ? n3249_o : 1'b0;
  /* decoder.vhd:1341:7  */
  assign n3271_o = opc_mnemonic_s == 6'b011101;
  /* decoder.vhd:1366:12  */
  assign n3272_o = ~clk_second_cycle_i;
  /* decoder.vhd:1368:27  */
  assign n3274_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1371:48  */
  assign n3275_o = opc_opcode_q[6];
  /* decoder.vhd:1368:11  */
  assign n3278_o = n3274_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1368:11  */
  assign n3281_o = n3274_o ? 1'b1 : 1'b0;
  assign n3282_o = opc_opcode_q[5];
  /* decoder.vhd:1366:9  */
  assign n3283_o = n3303_o ? n3275_o : n3282_o;
  /* decoder.vhd:1377:27  */
  assign n3285_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1377:37  */
  assign n3286_o = n3285_o & cnd_take_branch_i;
  /* decoder.vhd:1377:11  */
  assign n3292_o = n3286_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1377:11  */
  assign n3295_o = n3286_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1366:9  */
  assign n3297_o = n3272_o ? n3278_o : 1'b0;
  /* decoder.vhd:1366:9  */
  assign n3299_o = n3272_o ? 1'b0 : n3292_o;
  /* decoder.vhd:1366:9  */
  assign n3301_o = n3272_o ? n3281_o : 1'b0;
  /* decoder.vhd:1366:9  */
  assign n3303_o = n3272_o & n3274_o;
  /* decoder.vhd:1366:9  */
  assign n3305_o = n3272_o ? 1'b0 : n3295_o;
  /* decoder.vhd:1362:7  */
  assign n3307_o = opc_mnemonic_s == 6'b011110;
  /* decoder.vhd:1389:48  */
  assign n3309_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1389:31  */
  assign n3310_o = clk_second_cycle_i & n3309_o;
  /* decoder.vhd:1389:9  */
  assign n3313_o = n3310_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1384:7  */
  assign n3315_o = opc_mnemonic_s == 6'b011111;
  /* decoder.vhd:1399:28  */
  assign n3316_o = opc_opcode_q[3];
  /* decoder.vhd:1399:32  */
  assign n3317_o = ~n3316_o;
  /* decoder.vhd:1398:44  */
  assign n3319_o = 1'b0 | n3317_o;
  /* decoder.vhd:1398:13  */
  assign n3326_o = n3319_o ? 1'b1 : n2156_o;
  /* decoder.vhd:1398:13  */
  assign n3329_o = n3319_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1398:13  */
  assign n3332_o = n3319_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1397:11  */
  assign n3334_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1404:11  */
  assign n3339_o = clk_mstate_i == 3'b011;
  assign n3340_o = {n3339_o, n3334_o};
  /* decoder.vhd:1395:9  */
  always @*
    case (n3340_o)
      2'b10: n3343_o = 1'b1;
      2'b01: n3343_o = 1'b0;
      default: n3343_o = 1'b0;
    endcase
  /* decoder.vhd:1395:9  */
  always @*
    case (n3340_o)
      2'b10: n3346_o = 1'b1;
      2'b01: n3346_o = 1'b0;
      default: n3346_o = 1'b0;
    endcase
  /* decoder.vhd:1395:9  */
  always @*
    case (n3340_o)
      2'b10: n3347_o = n2156_o;
      2'b01: n3347_o = n3326_o;
      default: n3347_o = n2156_o;
    endcase
  /* decoder.vhd:1395:9  */
  always @*
    case (n3340_o)
      2'b10: n3350_o = 1'b1;
      2'b01: n3350_o = n3329_o;
      default: n3350_o = 1'b0;
    endcase
  /* decoder.vhd:1395:9  */
  always @*
    case (n3340_o)
      2'b10: n3352_o = 2'b01;
      2'b01: n3352_o = n3332_o;
      default: n3352_o = 2'b01;
    endcase
  /* decoder.vhd:1394:7  */
  assign n3354_o = opc_mnemonic_s == 6'b100001;
  /* decoder.vhd:1415:25  */
  assign n3356_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1415:9  */
  assign n3359_o = n3356_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1415:9  */
  assign n3362_o = n3356_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1415:9  */
  assign n3365_o = n3356_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1414:7  */
  assign n3367_o = opc_mnemonic_s == 6'b100000;
  /* decoder.vhd:1423:25  */
  assign n3369_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1423:9  */
  assign n3372_o = n3369_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1423:9  */
  assign n3375_o = n3369_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1423:9  */
  assign n3378_o = n3369_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1422:7  */
  assign n3380_o = opc_mnemonic_s == 6'b100010;
  /* decoder.vhd:1435:28  */
  assign n3381_o = opc_opcode_q[3];
  /* decoder.vhd:1435:32  */
  assign n3382_o = ~n3381_o;
  /* decoder.vhd:1434:44  */
  assign n3384_o = 1'b0 | n3382_o;
  /* decoder.vhd:1434:13  */
  assign n3391_o = n3384_o ? 1'b1 : n2156_o;
  /* decoder.vhd:1434:13  */
  assign n3394_o = n3384_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1434:13  */
  assign n3397_o = n3384_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1433:11  */
  assign n3399_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1440:11  */
  assign n3401_o = clk_mstate_i == 3'b100;
  assign n3402_o = {n3401_o, n3399_o};
  /* decoder.vhd:1431:9  */
  always @*
    case (n3402_o)
      2'b10: n3405_o = 1'b1;
      2'b01: n3405_o = 1'b0;
      default: n3405_o = 1'b0;
    endcase
  /* decoder.vhd:1431:9  */
  always @*
    case (n3402_o)
      2'b10: n3406_o = n2156_o;
      2'b01: n3406_o = n3391_o;
      default: n3406_o = n2156_o;
    endcase
  /* decoder.vhd:1431:9  */
  always @*
    case (n3402_o)
      2'b10: n3408_o = 1'b0;
      2'b01: n3408_o = n3394_o;
      default: n3408_o = 1'b0;
    endcase
  /* decoder.vhd:1431:9  */
  always @*
    case (n3402_o)
      2'b10: n3410_o = 2'b01;
      2'b01: n3410_o = n3397_o;
      default: n3410_o = 2'b01;
    endcase
  /* decoder.vhd:1431:9  */
  always @*
    case (n3402_o)
      2'b10: n3413_o = 1'b1;
      2'b01: n3413_o = 1'b0;
      default: n3413_o = 1'b0;
    endcase
  /* decoder.vhd:1430:7  */
  assign n3415_o = opc_mnemonic_s == 6'b100011;
  /* decoder.vhd:1454:12  */
  assign n3416_o = ~clk_second_cycle_i;
  /* decoder.vhd:1454:52  */
  assign n3418_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1454:35  */
  assign n3419_o = n3416_o & n3418_o;
  /* decoder.vhd:1456:26  */
  assign n3420_o = opc_opcode_q[3];
  /* decoder.vhd:1456:30  */
  assign n3421_o = ~n3420_o;
  /* decoder.vhd:1455:42  */
  assign n3423_o = 1'b0 | n3421_o;
  /* decoder.vhd:1454:9  */
  assign n3430_o = n3437_o ? 1'b1 : n2156_o;
  /* decoder.vhd:1455:11  */
  assign n3433_o = n3423_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1455:11  */
  assign n3436_o = n3423_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1454:9  */
  assign n3437_o = n3419_o & n3423_o;
  /* decoder.vhd:1454:9  */
  assign n3439_o = n3419_o ? n3433_o : 1'b0;
  /* decoder.vhd:1454:9  */
  assign n3441_o = n3419_o ? n3436_o : 2'b01;
  /* decoder.vhd:1463:48  */
  assign n3443_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1463:31  */
  assign n3444_o = clk_second_cycle_i & n3443_o;
  /* decoder.vhd:1463:9  */
  assign n3447_o = n3444_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1450:7  */
  assign n3449_o = opc_mnemonic_s == 6'b100100;
  /* decoder.vhd:1470:25  */
  assign n3451_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1470:9  */
  assign n3454_o = n3451_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1470:9  */
  assign n3457_o = n3451_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1468:7  */
  assign n3459_o = opc_mnemonic_s == 6'b111111;
  /* decoder.vhd:1478:25  */
  assign n3461_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1479:26  */
  assign n3462_o = opc_opcode_q[5];
  /* decoder.vhd:1479:11  */
  assign n3465_o = n3462_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1479:11  */
  assign n3468_o = n3462_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1479:11  */
  assign n3471_o = n3462_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1479:11  */
  assign n3474_o = n3462_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1478:9  */
  assign n3476_o = n3461_o ? n3465_o : 1'b0;
  /* decoder.vhd:1478:9  */
  assign n3478_o = n3461_o ? n3468_o : 1'b0;
  /* decoder.vhd:1478:9  */
  assign n3480_o = n3461_o ? n3471_o : 1'b0;
  /* decoder.vhd:1478:9  */
  assign n3482_o = n3461_o ? n3474_o : 1'b0;
  /* decoder.vhd:1477:7  */
  assign n3484_o = opc_mnemonic_s == 6'b100101;
  /* decoder.vhd:1492:12  */
  assign n3485_o = ~clk_second_cycle_i;
  /* decoder.vhd:1498:53  */
  assign n3487_o = opc_opcode_q[1:0];
  /* decoder.vhd:1500:32  */
  assign n3488_o = opc_opcode_q[7:4];
  /* decoder.vhd:1501:17  */
  assign n3491_o = n3488_o == 4'b1001;
  /* decoder.vhd:1503:17  */
  assign n3494_o = n3488_o == 4'b1000;
  /* decoder.vhd:1505:17  */
  assign n3497_o = n3488_o == 4'b0011;
  assign n3498_o = {n3497_o, n3494_o, n3491_o};
  assign n3499_o = n2158_o[3:2];
  assign n3500_o = n2159_o[3:2];
  /* decoder.vhd:622:5  */
  assign n3501_o = n2145_o ? n3499_o : n3500_o;
  /* decoder.vhd:1500:15  */
  always @*
    case (n3498_o)
      3'b100: n3502_o = 2'b01;
      3'b010: n3502_o = 2'b10;
      3'b001: n3502_o = 2'b11;
      default: n3502_o = n3501_o;
    endcase
  /* decoder.vhd:1495:13  */
  assign n3504_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1516:13  */
  assign n3506_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1522:13  */
  assign n3508_o = clk_mstate_i == 3'b100;
  assign n3509_o = {n3508_o, n3506_o, n3504_o};
  /* decoder.vhd:1493:11  */
  always @*
    case (n3509_o)
      3'b100: n3512_o = 1'b0;
      3'b010: n3512_o = 1'b1;
      3'b001: n3512_o = 1'b0;
      default: n3512_o = 1'b0;
    endcase
  /* decoder.vhd:1493:11  */
  always @*
    case (n3509_o)
      3'b100: n3516_o = 1'b0;
      3'b010: n3516_o = 1'b1;
      3'b001: n3516_o = 1'b1;
      default: n3516_o = 1'b0;
    endcase
  assign n3517_o = n2158_o[1:0];
  assign n3518_o = n2159_o[1:0];
  /* decoder.vhd:622:5  */
  assign n3519_o = n2145_o ? n3517_o : n3518_o;
  /* decoder.vhd:1493:11  */
  always @*
    case (n3509_o)
      3'b100: n3520_o = n3519_o;
      3'b010: n3520_o = n3519_o;
      3'b001: n3520_o = n3487_o;
      default: n3520_o = n3519_o;
    endcase
  assign n3521_o = n2158_o[3:2];
  assign n3522_o = n2159_o[3:2];
  /* decoder.vhd:622:5  */
  assign n3523_o = n2145_o ? n3521_o : n3522_o;
  /* decoder.vhd:1493:11  */
  always @*
    case (n3509_o)
      3'b100: n3524_o = n3523_o;
      3'b010: n3524_o = n3523_o;
      3'b001: n3524_o = n3502_o;
      default: n3524_o = n3523_o;
    endcase
  assign n3525_o = n2158_o[7:4];
  assign n3526_o = n2159_o[7:4];
  /* decoder.vhd:622:5  */
  assign n3527_o = n2145_o ? n3525_o : n3526_o;
  /* decoder.vhd:1493:11  */
  always @*
    case (n3509_o)
      3'b100: n3528_o = n3527_o;
      3'b010: n3528_o = n3527_o;
      3'b001: n3528_o = 4'b0000;
      default: n3528_o = n3527_o;
    endcase
  /* decoder.vhd:1493:11  */
  always @*
    case (n3509_o)
      3'b100: n3530_o = n2164_o;
      3'b010: n3530_o = n2164_o;
      3'b001: n3530_o = 1'b1;
      default: n3530_o = n2164_o;
    endcase
  /* decoder.vhd:1493:11  */
  always @*
    case (n3509_o)
      3'b100: n3534_o = 1'b1;
      3'b010: n3534_o = 1'b1;
      3'b001: n3534_o = 1'b0;
      default: n3534_o = 1'b0;
    endcase
  /* decoder.vhd:1532:27  */
  assign n3536_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1532:53  */
  assign n3538_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1532:37  */
  assign n3539_o = n3536_o | n3538_o;
  /* decoder.vhd:1532:11  */
  assign n3542_o = n3539_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1492:9  */
  assign n3544_o = n3485_o ? n3512_o : 1'b0;
  /* decoder.vhd:1492:9  */
  assign n3546_o = n3485_o ? n3516_o : 1'b0;
  assign n3547_o = {n3528_o, n3524_o, n3520_o};
  /* decoder.vhd:1492:9  */
  assign n3548_o = n3485_o ? n3547_o : n2160_o;
  /* decoder.vhd:1492:9  */
  assign n3549_o = n3485_o ? n3530_o : n2164_o;
  /* decoder.vhd:1492:9  */
  assign n3550_o = n3485_o ? n3534_o : n3542_o;
  /* decoder.vhd:1489:7  */
  assign n3552_o = opc_mnemonic_s == 6'b101101;
  /* decoder.vhd:1542:12  */
  assign n3553_o = ~clk_second_cycle_i;
  /* decoder.vhd:1548:53  */
  assign n3554_o = opc_opcode_q[1:0];
  /* decoder.vhd:1547:48  */
  assign n3556_o = {6'b000000, n3554_o};
  /* decoder.vhd:1545:13  */
  assign n3558_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1554:13  */
  assign n3561_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1561:13  */
  assign n3563_o = clk_mstate_i == 3'b100;
  assign n3564_o = {n3563_o, n3561_o, n3558_o};
  /* decoder.vhd:1543:11  */
  always @*
    case (n3564_o)
      3'b100: n3568_o = 1'b0;
      3'b010: n3568_o = 1'b1;
      3'b001: n3568_o = 1'b1;
      default: n3568_o = 1'b0;
    endcase
  assign n3569_o = n3556_o[3:0];
  assign n3570_o = n2158_o[3:0];
  assign n3571_o = n2159_o[3:0];
  /* decoder.vhd:622:5  */
  assign n3572_o = n2145_o ? n3570_o : n3571_o;
  /* decoder.vhd:1543:11  */
  always @*
    case (n3564_o)
      3'b100: n3573_o = n3572_o;
      3'b010: n3573_o = 4'b1111;
      3'b001: n3573_o = n3569_o;
      default: n3573_o = n3572_o;
    endcase
  assign n3574_o = n3556_o[7:4];
  assign n3575_o = n2158_o[7:4];
  assign n3576_o = n2159_o[7:4];
  /* decoder.vhd:622:5  */
  assign n3577_o = n2145_o ? n3575_o : n3576_o;
  /* decoder.vhd:1543:11  */
  always @*
    case (n3564_o)
      3'b100: n3578_o = n3577_o;
      3'b010: n3578_o = n3577_o;
      3'b001: n3578_o = n3574_o;
      default: n3578_o = n3577_o;
    endcase
  /* decoder.vhd:1543:11  */
  always @*
    case (n3564_o)
      3'b100: n3581_o = n2164_o;
      3'b010: n3581_o = 1'b1;
      3'b001: n3581_o = 1'b1;
      default: n3581_o = n2164_o;
    endcase
  /* decoder.vhd:1543:11  */
  always @*
    case (n3564_o)
      3'b100: n3585_o = 1'b1;
      3'b010: n3585_o = 1'b1;
      3'b001: n3585_o = 1'b0;
      default: n3585_o = 1'b0;
    endcase
  /* decoder.vhd:1572:13  */
  assign n3587_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1577:13  */
  assign n3589_o = clk_mstate_i == 3'b001;
  assign n3590_o = {n3589_o, n3587_o};
  /* decoder.vhd:1570:11  */
  always @*
    case (n3590_o)
      2'b10: n3593_o = 1'b1;
      2'b01: n3593_o = 1'b0;
      default: n3593_o = 1'b0;
    endcase
  /* decoder.vhd:1570:11  */
  always @*
    case (n3590_o)
      2'b10: n3596_o = 1'b1;
      2'b01: n3596_o = 1'b0;
      default: n3596_o = 1'b0;
    endcase
  /* decoder.vhd:1570:11  */
  always @*
    case (n3590_o)
      2'b10: n3599_o = 1'b1;
      2'b01: n3599_o = 1'b0;
      default: n3599_o = 1'b0;
    endcase
  /* decoder.vhd:1570:11  */
  always @*
    case (n3590_o)
      2'b10: n3603_o = 1'b1;
      2'b01: n3603_o = 1'b1;
      default: n3603_o = 1'b0;
    endcase
  /* decoder.vhd:1542:9  */
  assign n3605_o = n3553_o ? 1'b0 : n3593_o;
  /* decoder.vhd:1542:9  */
  assign n3607_o = n3553_o ? n3568_o : 1'b0;
  /* decoder.vhd:1542:9  */
  assign n3609_o = n3553_o ? 1'b0 : n3596_o;
  /* decoder.vhd:1542:9  */
  assign n3611_o = n3553_o ? 1'b0 : n3599_o;
  assign n3612_o = {n3578_o, n3573_o};
  /* decoder.vhd:1542:9  */
  assign n3613_o = n3553_o ? n3612_o : n2160_o;
  /* decoder.vhd:1542:9  */
  assign n3614_o = n3553_o ? n3581_o : n2164_o;
  /* decoder.vhd:1542:9  */
  assign n3615_o = n3553_o ? n3585_o : n3603_o;
  /* decoder.vhd:1539:7  */
  assign n3617_o = opc_mnemonic_s == 6'b100110;
  /* decoder.vhd:1594:12  */
  assign n3618_o = ~clk_second_cycle_i;
  /* decoder.vhd:1597:27  */
  assign n3620_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1599:28  */
  assign n3621_o = opc_opcode_q[6];
  /* decoder.vhd:1599:32  */
  assign n3622_o = ~n3621_o;
  /* decoder.vhd:1599:13  */
  assign n3625_o = n3622_o ? 2'b01 : 2'b10;
  /* decoder.vhd:1597:11  */
  assign n3628_o = n3620_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1597:11  */
  assign n3630_o = n3620_o ? n3625_o : 2'b00;
  /* decoder.vhd:1607:27  */
  assign n3632_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1607:11  */
  assign n3635_o = n3632_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1607:11  */
  assign n3638_o = n3632_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1594:9  */
  assign n3640_o = n3618_o ? 1'b0 : n3635_o;
  /* decoder.vhd:1594:9  */
  assign n3642_o = n3618_o ? n3628_o : 1'b0;
  /* decoder.vhd:1594:9  */
  assign n3644_o = n3618_o ? n3630_o : 2'b00;
  /* decoder.vhd:1594:9  */
  assign n3646_o = n3618_o ? 1'b0 : n3638_o;
  /* decoder.vhd:1591:7  */
  assign n3648_o = opc_mnemonic_s == 6'b100111;
  /* decoder.vhd:1621:24  */
  assign n3649_o = opc_opcode_q[4];
  /* decoder.vhd:1621:28  */
  assign n3650_o = ~n3649_o;
  /* decoder.vhd:1621:9  */
  assign n3653_o = n3650_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1621:9  */
  assign n3656_o = n3650_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1627:12  */
  assign n3657_o = ~clk_second_cycle_i;
  /* decoder.vhd:1631:13  */
  assign n3659_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1637:30  */
  assign n3660_o = opc_opcode_q[4];
  /* decoder.vhd:1637:15  */
  assign n3663_o = n3660_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1637:15  */
  assign n3666_o = n3660_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1636:13  */
  assign n3668_o = clk_mstate_i == 3'b100;
  assign n3669_o = {n3668_o, n3659_o};
  /* decoder.vhd:1629:11  */
  always @*
    case (n3669_o)
      2'b10: n3671_o = n3663_o;
      2'b01: n3671_o = 1'b0;
      default: n3671_o = 1'b0;
    endcase
  /* decoder.vhd:1629:11  */
  always @*
    case (n3669_o)
      2'b10: n3674_o = n3666_o;
      2'b01: n3674_o = 1'b1;
      default: n3674_o = 1'b0;
    endcase
  /* decoder.vhd:1629:11  */
  always @*
    case (n3669_o)
      2'b10: n3677_o = 1'b0;
      2'b01: n3677_o = 1'b1;
      default: n3677_o = 1'b0;
    endcase
  /* decoder.vhd:1647:27  */
  assign n3679_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1648:28  */
  assign n3680_o = opc_opcode_q[4];
  /* decoder.vhd:1648:32  */
  assign n3681_o = ~n3680_o;
  /* decoder.vhd:1648:13  */
  assign n3684_o = n3681_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1648:13  */
  assign n3687_o = n3681_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1648:13  */
  assign n3690_o = n3681_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1648:13  */
  assign n3693_o = n3681_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1647:11  */
  assign n3695_o = n3679_o ? n3684_o : 1'b0;
  /* decoder.vhd:1647:11  */
  assign n3697_o = n3679_o ? n3687_o : 1'b0;
  /* decoder.vhd:1647:11  */
  assign n3699_o = n3679_o ? n3690_o : 1'b0;
  /* decoder.vhd:1647:11  */
  assign n3701_o = n3679_o ? n3693_o : 1'b0;
  /* decoder.vhd:1627:9  */
  assign n3703_o = n3657_o ? 1'b0 : n3695_o;
  /* decoder.vhd:1627:9  */
  assign n3704_o = n3657_o ? n3671_o : n3697_o;
  /* decoder.vhd:1627:9  */
  assign n3705_o = n3657_o ? n3674_o : n3699_o;
  /* decoder.vhd:1627:9  */
  assign n3707_o = n3657_o ? n3677_o : 1'b0;
  /* decoder.vhd:1627:9  */
  assign n3709_o = n3657_o ? 1'b0 : n3701_o;
  /* decoder.vhd:1627:9  */
  assign n3712_o = n3657_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1618:7  */
  assign n3714_o = opc_mnemonic_s == 6'b101000;
  /* decoder.vhd:1663:7  */
  assign n3716_o = opc_mnemonic_s == 6'b101001;
  /* decoder.vhd:1672:28  */
  assign n3717_o = opc_opcode_q[3];
  /* decoder.vhd:1672:32  */
  assign n3718_o = ~n3717_o;
  /* decoder.vhd:1671:44  */
  assign n3720_o = 1'b0 | n3718_o;
  /* decoder.vhd:1671:13  */
  assign n3727_o = n3720_o ? 1'b1 : n2156_o;
  /* decoder.vhd:1671:13  */
  assign n3730_o = n3720_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1671:13  */
  assign n3733_o = n3720_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1670:11  */
  assign n3735_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1677:11  */
  assign n3740_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1681:11  */
  assign n3745_o = clk_mstate_i == 3'b100;
  assign n3746_o = {n3745_o, n3740_o, n3735_o};
  /* decoder.vhd:1668:9  */
  always @*
    case (n3746_o)
      3'b100: n3749_o = 1'b1;
      3'b010: n3749_o = 1'b0;
      3'b001: n3749_o = 1'b0;
      default: n3749_o = 1'b0;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3746_o)
      3'b100: n3752_o = 1'b0;
      3'b010: n3752_o = 1'b1;
      3'b001: n3752_o = 1'b0;
      default: n3752_o = 1'b0;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3746_o)
      3'b100: n3755_o = 1'b1;
      3'b010: n3755_o = 1'b0;
      3'b001: n3755_o = 1'b0;
      default: n3755_o = 1'b0;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3746_o)
      3'b100: n3756_o = n2156_o;
      3'b010: n3756_o = n2156_o;
      3'b001: n3756_o = n3727_o;
      default: n3756_o = n2156_o;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3746_o)
      3'b100: n3759_o = 1'b0;
      3'b010: n3759_o = 1'b1;
      3'b001: n3759_o = n3730_o;
      default: n3759_o = 1'b0;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3746_o)
      3'b100: n3762_o = 4'b0001;
      3'b010: n3762_o = 4'b1100;
      3'b001: n3762_o = 4'b1100;
      default: n3762_o = 4'b1100;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3746_o)
      3'b100: n3764_o = 2'b01;
      3'b010: n3764_o = 2'b01;
      3'b001: n3764_o = n3733_o;
      default: n3764_o = 2'b01;
    endcase
  /* decoder.vhd:1667:7  */
  assign n3766_o = opc_mnemonic_s == 6'b101010;
  /* decoder.vhd:1696:13  */
  assign n3768_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1700:13  */
  assign n3773_o = clk_mstate_i == 3'b010;
  assign n3774_o = {n3773_o, n3768_o};
  /* decoder.vhd:1694:11  */
  always @*
    case (n3774_o)
      2'b10: n3777_o = 1'b1;
      2'b01: n3777_o = 1'b0;
      default: n3777_o = 1'b0;
    endcase
  /* decoder.vhd:1694:11  */
  always @*
    case (n3774_o)
      2'b10: n3780_o = 1'b0;
      2'b01: n3780_o = 1'b1;
      default: n3780_o = 1'b0;
    endcase
  /* decoder.vhd:1694:11  */
  always @*
    case (n3774_o)
      2'b10: n3783_o = 1'b1;
      2'b01: n3783_o = 1'b0;
      default: n3783_o = 1'b0;
    endcase
  /* decoder.vhd:1694:11  */
  always @*
    case (n3774_o)
      2'b10: n3786_o = 4'b0001;
      2'b01: n3786_o = 4'b1100;
      default: n3786_o = 4'b1100;
    endcase
  /* decoder.vhd:1693:9  */
  assign n3788_o = clk_second_cycle_i ? n3777_o : 1'b0;
  /* decoder.vhd:1693:9  */
  assign n3790_o = clk_second_cycle_i ? n3780_o : 1'b0;
  /* decoder.vhd:1693:9  */
  assign n3792_o = clk_second_cycle_i ? n3783_o : 1'b0;
  /* decoder.vhd:1693:9  */
  assign n3794_o = clk_second_cycle_i ? n3786_o : 4'b1100;
  /* decoder.vhd:1690:7  */
  assign n3796_o = opc_mnemonic_s == 6'b101011;
  /* decoder.vhd:1714:12  */
  assign n3797_o = ~clk_second_cycle_i;
  /* decoder.vhd:1716:27  */
  assign n3799_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:1717:28  */
  assign n3800_o = opc_opcode_q[1:0];
  /* decoder.vhd:1717:41  */
  assign n3802_o = n3800_o == 2'b00;
  /* decoder.vhd:1719:31  */
  assign n3803_o = opc_opcode_q[1];
  /* decoder.vhd:1719:35  */
  assign n3804_o = ~n3803_o;
  /* decoder.vhd:1719:13  */
  assign n3807_o = n3804_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1719:13  */
  assign n3810_o = n3804_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1719:13  */
  assign n3813_o = n3804_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1719:13  */
  assign n3816_o = n3804_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1717:13  */
  assign n3818_o = n3802_o ? 1'b0 : n3807_o;
  /* decoder.vhd:1717:13  */
  assign n3820_o = n3802_o ? 1'b0 : n3810_o;
  /* decoder.vhd:1717:13  */
  assign n3822_o = n3802_o ? 1'b0 : n3813_o;
  /* decoder.vhd:1717:13  */
  assign n3824_o = n3802_o ? 1'b0 : n3816_o;
  /* decoder.vhd:1717:13  */
  assign n3827_o = n3802_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3830_o = n3799_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3832_o = n3799_o ? n3818_o : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3834_o = n3799_o ? n3820_o : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3836_o = n3799_o ? n3822_o : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3838_o = n3799_o ? n3824_o : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3840_o = n3799_o ? n3827_o : 1'b0;
  /* decoder.vhd:1734:13  */
  assign n3842_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1739:13  */
  assign n3844_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1748:30  */
  assign n3845_o = opc_opcode_q[1:0];
  /* decoder.vhd:1748:43  */
  assign n3847_o = n3845_o == 2'b00;
  /* decoder.vhd:1750:33  */
  assign n3848_o = opc_opcode_q[1];
  /* decoder.vhd:1750:37  */
  assign n3849_o = ~n3848_o;
  /* decoder.vhd:1750:15  */
  assign n3852_o = n3849_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1750:15  */
  assign n3855_o = n3849_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1748:15  */
  assign n3858_o = n3847_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1748:15  */
  assign n3860_o = n3847_o ? 1'b0 : n3852_o;
  /* decoder.vhd:1748:15  */
  assign n3862_o = n3847_o ? 1'b0 : n3855_o;
  /* decoder.vhd:1744:13  */
  assign n3864_o = clk_mstate_i == 3'b010;
  assign n3865_o = {n3864_o, n3844_o, n3842_o};
  /* decoder.vhd:1731:11  */
  always @*
    case (n3865_o)
      3'b100: n3869_o = 1'b0;
      3'b010: n3869_o = 1'b1;
      3'b001: n3869_o = 1'b1;
      default: n3869_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3865_o)
      3'b100: n3873_o = 1'b1;
      3'b010: n3873_o = 1'b1;
      3'b001: n3873_o = 1'b0;
      default: n3873_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3865_o)
      3'b100: n3875_o = n3858_o;
      3'b010: n3875_o = 1'b0;
      3'b001: n3875_o = 1'b0;
      default: n3875_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3865_o)
      3'b100: n3877_o = n3860_o;
      3'b010: n3877_o = 1'b0;
      3'b001: n3877_o = 1'b0;
      default: n3877_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3865_o)
      3'b100: n3879_o = n3862_o;
      3'b010: n3879_o = 1'b0;
      3'b001: n3879_o = 1'b0;
      default: n3879_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3865_o)
      3'b100: n3882_o = 4'b0001;
      3'b010: n3882_o = 4'b1100;
      3'b001: n3882_o = 4'b1100;
      default: n3882_o = 4'b1100;
    endcase
  /* decoder.vhd:1714:9  */
  assign n3884_o = n3797_o ? 1'b0 : n3869_o;
  /* decoder.vhd:1714:9  */
  assign n3886_o = n3797_o ? n3830_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3888_o = n3797_o ? 1'b0 : n3873_o;
  /* decoder.vhd:1714:9  */
  assign n3890_o = n3797_o ? 1'b0 : n3875_o;
  /* decoder.vhd:1714:9  */
  assign n3892_o = n3797_o ? 1'b0 : n3877_o;
  /* decoder.vhd:1714:9  */
  assign n3894_o = n3797_o ? n3832_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3896_o = n3797_o ? 1'b0 : n3879_o;
  /* decoder.vhd:1714:9  */
  assign n3898_o = n3797_o ? n3834_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3900_o = n3797_o ? 4'b1100 : n3882_o;
  /* decoder.vhd:1714:9  */
  assign n3902_o = n3797_o ? n3836_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3904_o = n3797_o ? n3838_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3906_o = n3797_o ? n3840_o : 1'b0;
  /* decoder.vhd:1711:7  */
  assign n3908_o = opc_mnemonic_s == 6'b101100;
  /* decoder.vhd:1766:25  */
  assign n3910_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1766:9  */
  assign n3913_o = n3910_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1766:9  */
  assign n3916_o = n3910_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1764:7  */
  assign n3918_o = opc_mnemonic_s == 6'b111011;
  /* decoder.vhd:1774:24  */
  assign n3919_o = opc_opcode_q[4];
  /* decoder.vhd:1774:28  */
  assign n3920_o = ~n3919_o;
  /* decoder.vhd:1774:9  */
  assign n3923_o = n3920_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1779:12  */
  assign n3924_o = ~clk_second_cycle_i;
  /* decoder.vhd:1779:52  */
  assign n3926_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1779:35  */
  assign n3927_o = n3924_o & n3926_o;
  /* decoder.vhd:1782:26  */
  assign n3928_o = opc_opcode_q[4];
  /* decoder.vhd:1783:28  */
  assign n3929_o = opc_opcode_q[1];
  /* decoder.vhd:1783:32  */
  assign n3930_o = ~n3929_o;
  /* decoder.vhd:1783:13  */
  assign n3933_o = n3930_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1783:13  */
  assign n3936_o = n3930_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1782:11  */
  assign n3939_o = n3928_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1782:11  */
  assign n3941_o = n3928_o ? n3933_o : 1'b0;
  /* decoder.vhd:1782:11  */
  assign n3943_o = n3928_o ? n3936_o : 1'b0;
  /* decoder.vhd:1779:9  */
  assign n3946_o = n3927_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1779:9  */
  assign n3948_o = n3927_o ? n3939_o : 1'b0;
  /* decoder.vhd:1779:9  */
  assign n3950_o = n3927_o ? n3941_o : 1'b0;
  /* decoder.vhd:1779:9  */
  assign n3952_o = n3927_o ? n3943_o : 1'b0;
  /* decoder.vhd:1773:7  */
  assign n3954_o = opc_mnemonic_s == 6'b101110;
  /* decoder.vhd:1798:12  */
  assign n3955_o = ~clk_second_cycle_i;
  /* decoder.vhd:1801:13  */
  assign n3957_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1805:13  */
  assign n3959_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1812:13  */
  assign n3961_o = clk_mstate_i == 3'b100;
  assign n3962_o = {n3961_o, n3959_o, n3957_o};
  /* decoder.vhd:1799:11  */
  always @*
    case (n3962_o)
      3'b100: n3965_o = 1'b1;
      3'b010: n3965_o = 1'b1;
      3'b001: n3965_o = n2156_o;
      default: n3965_o = n2156_o;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3962_o)
      3'b100: n3968_o = 1'b1;
      3'b010: n3968_o = 1'b0;
      3'b001: n3968_o = 1'b0;
      default: n3968_o = 1'b0;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3962_o)
      3'b100: n3971_o = 1'b1;
      3'b010: n3971_o = 1'b0;
      3'b001: n3971_o = 1'b0;
      default: n3971_o = 1'b0;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3962_o)
      3'b100: n3974_o = 1'b0;
      3'b010: n3974_o = 1'b1;
      3'b001: n3974_o = 1'b0;
      default: n3974_o = 1'b0;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3962_o)
      3'b100: n3978_o = 2'b11;
      3'b010: n3978_o = 2'b10;
      3'b001: n3978_o = 2'b01;
      default: n3978_o = 2'b01;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3962_o)
      3'b100: n3981_o = 1'b0;
      3'b010: n3981_o = 1'b0;
      3'b001: n3981_o = 1'b1;
      default: n3981_o = 1'b0;
    endcase
  /* decoder.vhd:1829:30  */
  assign n3982_o = opc_opcode_q[4];
  /* decoder.vhd:1829:15  */
  assign n3985_o = n3982_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1829:15  */
  assign n3988_o = n3982_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1826:13  */
  assign n3990_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1834:13  */
  assign n3992_o = clk_mstate_i == 3'b001;
  assign n3993_o = {n3992_o, n3990_o};
  /* decoder.vhd:1824:11  */
  always @*
    case (n3993_o)
      2'b10: n3996_o = 1'b0;
      2'b01: n3996_o = 1'b1;
      default: n3996_o = 1'b0;
    endcase
  /* decoder.vhd:1824:11  */
  always @*
    case (n3993_o)
      2'b10: n3999_o = 1'b0;
      2'b01: n3999_o = 1'b1;
      default: n3999_o = 1'b0;
    endcase
  /* decoder.vhd:1824:11  */
  always @*
    case (n3993_o)
      2'b10: n4001_o = 1'b0;
      2'b01: n4001_o = n3985_o;
      default: n4001_o = 1'b0;
    endcase
  /* decoder.vhd:1824:11  */
  always @*
    case (n3993_o)
      2'b10: n4004_o = 1'b1;
      2'b01: n4004_o = 1'b0;
      default: n4004_o = 1'b0;
    endcase
  /* decoder.vhd:1824:11  */
  always @*
    case (n3993_o)
      2'b10: n4006_o = 1'b0;
      2'b01: n4006_o = n3988_o;
      default: n4006_o = 1'b0;
    endcase
  /* decoder.vhd:1798:9  */
  assign n4007_o = n3955_o ? n3965_o : n2156_o;
  /* decoder.vhd:1798:9  */
  assign n4008_o = n3955_o ? n3968_o : n3996_o;
  /* decoder.vhd:1798:9  */
  assign n4010_o = n3955_o ? n3971_o : 1'b0;
  /* decoder.vhd:1798:9  */
  assign n4012_o = n3955_o ? 1'b0 : n3999_o;
  /* decoder.vhd:1798:9  */
  assign n4014_o = n3955_o ? n3974_o : 1'b0;
  /* decoder.vhd:1798:9  */
  assign n4016_o = n3955_o ? 1'b0 : n4001_o;
  /* decoder.vhd:1798:9  */
  assign n4018_o = n3955_o ? n3978_o : 2'b01;
  /* decoder.vhd:1798:9  */
  assign n4020_o = n3955_o ? n3981_o : 1'b0;
  /* decoder.vhd:1798:9  */
  assign n4022_o = n3955_o ? 1'b0 : n4004_o;
  /* decoder.vhd:1798:9  */
  assign n4024_o = n3955_o ? 1'b0 : n4006_o;
  /* decoder.vhd:1797:7  */
  assign n4026_o = opc_mnemonic_s == 6'b101111;
  /* decoder.vhd:1846:25  */
  assign n4028_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1851:26  */
  assign n4029_o = opc_opcode_q[4];
  /* decoder.vhd:1851:11  */
  assign n4032_o = n4029_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1851:11  */
  assign n4034_o = n4029_o ? alu_carry_i : 1'b0;
  /* decoder.vhd:1851:11  */
  assign n4037_o = n4029_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n4040_o = n4028_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n4043_o = n4028_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n4046_o = n4028_o ? 4'b0101 : 4'b1100;
  /* decoder.vhd:1846:9  */
  assign n4048_o = n4028_o ? n4032_o : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n4050_o = n4028_o ? n4034_o : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n4052_o = n4028_o ? n4037_o : 1'b0;
  /* decoder.vhd:1845:7  */
  assign n4054_o = opc_mnemonic_s == 6'b110000;
  /* decoder.vhd:1860:25  */
  assign n4056_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1865:26  */
  assign n4057_o = opc_opcode_q[4];
  /* decoder.vhd:1865:30  */
  assign n4058_o = ~n4057_o;
  /* decoder.vhd:1865:11  */
  assign n4061_o = n4058_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1865:11  */
  assign n4063_o = n4058_o ? alu_carry_i : 1'b0;
  /* decoder.vhd:1865:11  */
  assign n4066_o = n4058_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n4069_o = n4056_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n4072_o = n4056_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n4075_o = n4056_o ? 4'b0110 : 4'b1100;
  /* decoder.vhd:1860:9  */
  assign n4077_o = n4056_o ? n4061_o : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n4079_o = n4056_o ? n4063_o : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n4081_o = n4056_o ? n4066_o : 1'b0;
  /* decoder.vhd:1859:7  */
  assign n4083_o = opc_mnemonic_s == 6'b110001;
  /* decoder.vhd:1874:25  */
  assign n4085_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1875:26  */
  assign n4086_o = opc_opcode_q[4];
  /* decoder.vhd:1875:11  */
  assign n4089_o = n4086_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1875:11  */
  assign n4092_o = n4086_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1874:9  */
  assign n4094_o = n4085_o ? n4089_o : 1'b0;
  /* decoder.vhd:1874:9  */
  assign n4096_o = n4085_o ? n4092_o : 1'b0;
  /* decoder.vhd:1873:7  */
  assign n4098_o = opc_mnemonic_s == 6'b110010;
  /* decoder.vhd:1884:25  */
  assign n4100_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1885:45  */
  assign n4101_o = opc_opcode_q[4];
  /* decoder.vhd:1884:9  */
  assign n4103_o = n4100_o ? n4101_o : 1'b0;
  /* decoder.vhd:1884:9  */
  assign n4106_o = n4100_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1883:7  */
  assign n4108_o = opc_mnemonic_s == 6'b110011;
  /* decoder.vhd:1891:25  */
  assign n4110_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1891:9  */
  assign n4113_o = n4110_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1890:7  */
  assign n4115_o = opc_mnemonic_s == 6'b110100;
  /* decoder.vhd:1897:25  */
  assign n4117_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1898:26  */
  assign n4118_o = opc_opcode_q[4];
  /* decoder.vhd:1898:11  */
  assign n4121_o = n4118_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1898:11  */
  assign n4124_o = n4118_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1897:9  */
  assign n4126_o = n4117_o ? n4121_o : 1'b0;
  /* decoder.vhd:1897:9  */
  assign n4128_o = n4117_o ? n4124_o : 1'b0;
  /* decoder.vhd:1896:7  */
  assign n4130_o = opc_mnemonic_s == 6'b110101;
  /* decoder.vhd:1909:25  */
  assign n4132_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1909:9  */
  assign n4135_o = n4132_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1909:9  */
  assign n4138_o = n4132_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1906:7  */
  assign n4140_o = opc_mnemonic_s == 6'b110110;
  /* decoder.vhd:1920:28  */
  assign n4141_o = opc_opcode_q[3];
  /* decoder.vhd:1920:32  */
  assign n4142_o = ~n4141_o;
  /* decoder.vhd:1919:44  */
  assign n4144_o = 1'b0 | n4142_o;
  /* decoder.vhd:1919:13  */
  assign n4151_o = n4144_o ? 1'b1 : n2156_o;
  /* decoder.vhd:1919:13  */
  assign n4154_o = n4144_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1919:13  */
  assign n4157_o = n4144_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1918:11  */
  assign n4159_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1930:28  */
  assign n4160_o = opc_opcode_q[4];
  /* decoder.vhd:1930:13  */
  assign n4163_o = n4160_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1926:11  */
  assign n4165_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1940:28  */
  assign n4166_o = opc_opcode_q[4];
  /* decoder.vhd:1940:13  */
  assign n4169_o = n4166_o ? 4'b1011 : 4'b1100;
  /* decoder.vhd:1937:11  */
  assign n4171_o = clk_mstate_i == 3'b100;
  assign n4172_o = {n4171_o, n4165_o, n4159_o};
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4175_o = 1'b0;
      3'b010: n4175_o = 1'b1;
      3'b001: n4175_o = 1'b0;
      default: n4175_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4178_o = 1'b0;
      3'b010: n4178_o = 1'b1;
      3'b001: n4178_o = 1'b0;
      default: n4178_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4181_o = 1'b1;
      3'b010: n4181_o = 1'b0;
      3'b001: n4181_o = 1'b0;
      default: n4181_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4182_o = n2156_o;
      3'b010: n4182_o = n2156_o;
      3'b001: n4182_o = n4151_o;
      default: n4182_o = n2156_o;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4185_o = 1'b0;
      3'b010: n4185_o = 1'b1;
      3'b001: n4185_o = n4154_o;
      default: n4185_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4187_o = n4169_o;
      3'b010: n4187_o = 4'b1100;
      3'b001: n4187_o = 4'b1100;
      default: n4187_o = 4'b1100;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4189_o = 1'b0;
      3'b010: n4189_o = n4163_o;
      3'b001: n4189_o = 1'b0;
      default: n4189_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4191_o = 2'b01;
      3'b010: n4191_o = 2'b01;
      3'b001: n4191_o = n4157_o;
      default: n4191_o = 2'b01;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4172_o)
      3'b100: n4194_o = 1'b1;
      3'b010: n4194_o = 1'b0;
      3'b001: n4194_o = 1'b0;
      default: n4194_o = 1'b0;
    endcase
  /* decoder.vhd:1915:7  */
  assign n4196_o = opc_mnemonic_s == 6'b110111;
  /* decoder.vhd:1957:28  */
  assign n4197_o = opc_opcode_q[3];
  /* decoder.vhd:1957:32  */
  assign n4198_o = ~n4197_o;
  /* decoder.vhd:1956:44  */
  assign n4200_o = 1'b0 | n4198_o;
  /* decoder.vhd:1956:13  */
  assign n4207_o = n4200_o ? 1'b1 : n2156_o;
  /* decoder.vhd:1956:13  */
  assign n4210_o = n4200_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1956:13  */
  assign n4213_o = n4200_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1955:11  */
  assign n4215_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1962:11  */
  assign n4220_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1966:11  */
  assign n4225_o = clk_mstate_i == 3'b100;
  assign n4226_o = {n4225_o, n4220_o, n4215_o};
  /* decoder.vhd:1953:9  */
  always @*
    case (n4226_o)
      3'b100: n4229_o = 1'b1;
      3'b010: n4229_o = 1'b0;
      3'b001: n4229_o = 1'b0;
      default: n4229_o = 1'b0;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4226_o)
      3'b100: n4232_o = 1'b0;
      3'b010: n4232_o = 1'b1;
      3'b001: n4232_o = 1'b0;
      default: n4232_o = 1'b0;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4226_o)
      3'b100: n4235_o = 1'b1;
      3'b010: n4235_o = 1'b0;
      3'b001: n4235_o = 1'b0;
      default: n4235_o = 1'b0;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4226_o)
      3'b100: n4236_o = n2156_o;
      3'b010: n4236_o = n2156_o;
      3'b001: n4236_o = n4207_o;
      default: n4236_o = n2156_o;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4226_o)
      3'b100: n4239_o = 1'b0;
      3'b010: n4239_o = 1'b1;
      3'b001: n4239_o = n4210_o;
      default: n4239_o = 1'b0;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4226_o)
      3'b100: n4242_o = 4'b0010;
      3'b010: n4242_o = 4'b1100;
      3'b001: n4242_o = 4'b1100;
      default: n4242_o = 4'b1100;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4226_o)
      3'b100: n4244_o = 2'b01;
      3'b010: n4244_o = 2'b01;
      3'b001: n4244_o = n4213_o;
      default: n4244_o = 2'b01;
    endcase
  /* decoder.vhd:1952:7  */
  assign n4246_o = opc_mnemonic_s == 6'b111000;
  /* decoder.vhd:1981:13  */
  assign n4248_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1985:13  */
  assign n4253_o = clk_mstate_i == 3'b010;
  assign n4254_o = {n4253_o, n4248_o};
  /* decoder.vhd:1979:11  */
  always @*
    case (n4254_o)
      2'b10: n4257_o = 1'b1;
      2'b01: n4257_o = 1'b0;
      default: n4257_o = 1'b0;
    endcase
  /* decoder.vhd:1979:11  */
  always @*
    case (n4254_o)
      2'b10: n4260_o = 1'b0;
      2'b01: n4260_o = 1'b1;
      default: n4260_o = 1'b0;
    endcase
  /* decoder.vhd:1979:11  */
  always @*
    case (n4254_o)
      2'b10: n4263_o = 1'b1;
      2'b01: n4263_o = 1'b0;
      default: n4263_o = 1'b0;
    endcase
  /* decoder.vhd:1979:11  */
  always @*
    case (n4254_o)
      2'b10: n4266_o = 4'b0010;
      2'b01: n4266_o = 4'b1100;
      default: n4266_o = 4'b1100;
    endcase
  /* decoder.vhd:1978:9  */
  assign n4268_o = clk_second_cycle_i ? n4257_o : 1'b0;
  /* decoder.vhd:1978:9  */
  assign n4270_o = clk_second_cycle_i ? n4260_o : 1'b0;
  /* decoder.vhd:1978:9  */
  assign n4272_o = clk_second_cycle_i ? n4263_o : 1'b0;
  /* decoder.vhd:1978:9  */
  assign n4274_o = clk_second_cycle_i ? n4266_o : 4'b1100;
  /* decoder.vhd:1975:7  */
  assign n4276_o = opc_mnemonic_s == 6'b111001;
  assign n4277_o = {n4276_o, n4246_o, n4196_o, n4140_o, n4130_o, n4115_o, n4108_o, n4098_o, n4083_o, n4054_o, n4026_o, n3954_o, n3918_o, n3908_o, n3796_o, n3766_o, n3716_o, n3714_o, n3648_o, n3617_o, n3552_o, n3484_o, n3459_o, n3449_o, n3415_o, n3380_o, n3367_o, n3354_o, n3315_o, n3307_o, n3271_o, n3240_o, n3204_o, n3178_o, n3152_o, n3126_o, n3099_o, n3068_o, n3034_o, n3003_o, n2972_o, n2911_o, n2900_o, n2890_o, n2870_o, n2863_o, n2847_o, n2783_o, n2768_o, n2753_o, n2717_o, n2671_o, n2650_o, n2640_o, n2627_o, n2611_o, n2604_o, n2591_o, n2473_o, n2361_o, n2331_o, n2281_o, n2229_o};
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4279_o = n4268_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4279_o = n4229_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4279_o = n4175_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4279_o = n4135_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4279_o = n4069_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4279_o = n4040_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4279_o = n3788_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4279_o = n3749_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4279_o = n3703_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4279_o = n3640_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4279_o = n3605_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4279_o = n3476_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4279_o = n3359_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4279_o = n3343_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4279_o = n3313_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4279_o = n2955_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4279_o = n2906_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4279_o = n2895_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4279_o = n2884_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4279_o = n2739_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4279_o = n2693_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4279_o = n2632_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4279_o = n2596_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4279_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4279_o = n2353_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4279_o = n2314_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4279_o = n2265_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4279_o = n2202_o;
      default: n4279_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4282_o = n3884_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4282_o = n2957_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4282_o = n2827_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4282_o = n2741_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4282_o = n2695_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4282_o = n2449_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4282_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4282_o = 1'b0;
      default: n4282_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4285_o = n4270_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4285_o = n4232_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4285_o = n4178_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4285_o = n3886_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4285_o = n3790_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4285_o = n3752_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4285_o = n3346_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4285_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4285_o = n2451_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4285_o = n2355_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4285_o = n2317_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4285_o = n2267_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4285_o = n2205_o;
      default: n4285_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4288_o = n4272_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4288_o = n4235_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4288_o = n4181_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4288_o = n4138_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4288_o = n4072_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4288_o = n4043_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4288_o = n3946_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4288_o = n3913_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4288_o = n3888_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4288_o = n3792_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4288_o = n3755_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4288_o = n3704_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4288_o = n3642_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4288_o = n3544_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4288_o = n3478_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4288_o = n3454_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4288_o = n3405_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4288_o = n3372_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4288_o = n3297_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4288_o = n3118_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4288_o = n2995_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4288_o = n2960_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4288_o = n2829_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4288_o = n2744_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4288_o = n2698_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4288_o = n2635_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4288_o = n2599_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4288_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4288_o = n2453_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4288_o = n2357_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4288_o = n2320_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4288_o = n2269_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4288_o = n2208_o;
      default: n4288_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4291_o = n3948_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4291_o = n3916_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4291_o = n3890_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4291_o = n3705_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4291_o = n2455_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4291_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4291_o = 1'b0;
      default: n4291_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4294_o = n2562_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4294_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4294_o = 1'b0;
      default: n4294_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4297_o = n2859_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4297_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4297_o = 1'b0;
      default: n4297_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4300_o = n2861_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4300_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4300_o = 1'b0;
      default: n4300_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4303_o = n3457_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4303_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4303_o = 1'b0;
      default: n4303_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4305_o = n4236_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4305_o = n4182_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4305_o = n4007_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4305_o = n3756_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4305_o = n3430_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4305_o = n3406_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4305_o = n3347_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4305_o = n2961_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4305_o = n2563_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4305_o = n2321_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4305_o = n2156_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4305_o = n2209_o;
      default: n4305_o = n2156_o;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4307_o = n4239_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4307_o = n4185_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4307_o = n4008_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4307_o = n3759_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4307_o = n3707_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4307_o = n3439_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4307_o = n3408_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4307_o = n3350_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4307_o = n2963_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4307_o = n2831_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4307_o = n2746_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4307_o = n2324_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4307_o = n2212_o;
      default: n4307_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4310_o = n3950_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4310_o = n3892_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4310_o = n2457_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4310_o = 1'b0;
      default: n4310_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4313_o = n3894_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4313_o = n2886_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4313_o = n2459_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4313_o = 1'b0;
      default: n4313_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4316_o = n3952_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4316_o = n3896_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4316_o = n2461_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4316_o = 1'b0;
      default: n4316_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4319_o = n3607_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4319_o = n3546_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4319_o = 1'b0;
      default: n4319_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4322_o = n3898_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4322_o = n3609_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4322_o = n2888_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4322_o = n2463_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4322_o = 1'b0;
      default: n4322_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4325_o = n3611_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4325_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4325_o = 1'b0;
      default: n4325_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4328_o = n4010_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4328_o = n3299_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4328_o = n3263_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4328_o = n3232_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4328_o = n3198_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4328_o = n3172_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4328_o = n3146_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4328_o = n3120_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4328_o = n3091_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4328_o = n3060_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4328_o = n3026_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4328_o = n2997_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4328_o = n2833_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4328_o = n2565_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4328_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4328_o = 1'b0;
      default: n4328_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4331_o = n2567_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4331_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4331_o = 1'b0;
      default: n4331_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4334_o = n4012_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4334_o = n3093_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4334_o = n2569_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4334_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4334_o = 1'b0;
      default: n4334_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4337_o = n2571_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4337_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4337_o = 1'b0;
      default: n4337_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4340_o = n3362_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4340_o = n2573_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4340_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4340_o = 1'b0;
      default: n4340_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4343_o = n4014_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4343_o = n3365_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4343_o = n2575_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4343_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4343_o = 1'b0;
      default: n4343_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4346_o = n4016_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4346_o = n3375_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4346_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4346_o = 1'b0;
      default: n4346_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4349_o = n3378_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4349_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4349_o = 1'b0;
      default: n4349_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4353_o = n4274_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4353_o = n4242_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4353_o = n4187_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4353_o = 4'b0111;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4353_o = n4075_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4353_o = n4046_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4353_o = n3900_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4353_o = n3794_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4353_o = n3762_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4353_o = n2966_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4353_o = n2835_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4353_o = n2749_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4353_o = n2700_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4353_o = n2638_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4353_o = n2602_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4353_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4353_o = n2465_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4353_o = n2359_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4353_o = n2327_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4353_o = n2271_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4353_o = n2215_o;
      default: n4353_o = 4'b1100;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4356_o = n4077_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4356_o = n4048_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4356_o = n2273_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4356_o = n2217_o;
      default: n4356_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4359_o = n2704_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4359_o = 1'b0;
      default: n4359_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4362_o = n4189_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4362_o = 1'b0;
      default: n4362_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4365_o = n2707_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4365_o = 1'b0;
      default: n4365_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4368_o = n2710_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4368_o = 1'b0;
      default: n4368_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4372_o = 1'b1;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4372_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4372_o = 1'b0;
      default: n4372_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4377_o = 1'b1;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4377_o = 1'b1;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4377_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4377_o = 1'b0;
      default: n4377_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4381_o = n3653_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4381_o = 1'b1;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4381_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4381_o = 1'b0;
      default: n4381_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4384_o = n3923_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4384_o = n3656_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4384_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4384_o = 1'b0;
      default: n4384_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4387_o = n3301_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4387_o = n3265_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4387_o = n3234_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4387_o = n3200_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4387_o = n3174_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4387_o = n3148_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4387_o = n3062_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4387_o = n3028_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4387_o = n2999_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4387_o = n2837_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4387_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4387_o = 1'b0;
      default: n4387_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4397_o = 4'b0001;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4397_o = 4'b1000;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4397_o = n3209_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4397_o = 4'b1010;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4397_o = 4'b1001;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4397_o = 4'b0101;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4397_o = n3064_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4397_o = 4'b0010;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4397_o = n2839_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4397_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4397_o = 4'b0000;
      default: n4397_o = 4'b0000;
    endcase
  assign n4399_o = opc_opcode_q[5];
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4400_o = n3283_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4400_o = n3218_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4400_o = n3012_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4400_o = n2841_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4400_o = n4399_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4400_o = n4399_o;
      default: n4400_o = n4399_o;
    endcase
  assign n4401_o = opc_opcode_q[7:6];
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4403_o = n4244_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4403_o = n4191_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4403_o = n4018_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4403_o = n3764_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4403_o = n3441_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4403_o = n3410_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4403_o = n3352_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4403_o = n2968_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4403_o = n2577_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4403_o = n2329_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4403_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4403_o = n2219_o;
      default: n4403_o = 2'b01;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4406_o = n3902_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4406_o = n2467_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4406_o = 1'b0;
      default: n4406_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4409_o = n3904_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4409_o = n2469_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4409_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4409_o = 1'b0;
      default: n4409_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4412_o = n3644_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4412_o = n3122_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4412_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4412_o = 2'b00;
      default: n4412_o = 2'b00;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4415_o = n4103_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4415_o = n4079_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4415_o = n4050_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4415_o = n2712_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4415_o = n2665_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4415_o = n2645_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4415_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4415_o = n2275_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4415_o = n2221_o;
      default: n4415_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4418_o = n2579_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4418_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4418_o = 1'b0;
      default: n4418_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4421_o = n4020_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4421_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4421_o = 1'b0;
      default: n4421_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4424_o = n4081_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4424_o = n4052_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4424_o = n2715_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4424_o = n2648_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4424_o = n2609_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4424_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4424_o = n2277_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4424_o = n2224_o;
      default: n4424_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4427_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4427_o = n2279_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4427_o = n2227_o;
      default: n4427_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4430_o = n2667_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4430_o = n2623_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4430_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4430_o = 1'b0;
      default: n4430_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4433_o = n4106_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4433_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4433_o = 1'b0;
      default: n4433_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4436_o = n3480_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4436_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4436_o = 1'b0;
      default: n4436_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4439_o = n3482_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4439_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4439_o = 1'b0;
      default: n4439_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4442_o = n4126_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4442_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4442_o = 1'b0;
      default: n4442_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4445_o = n4128_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4445_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4445_o = 1'b0;
      default: n4445_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4448_o = n4113_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4448_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4448_o = 1'b0;
      default: n4448_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4473_o = 1'b1;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4473_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4473_o = 1'b1;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4473_o = 1'b0;
      default: n4473_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4476_o = n3646_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4476_o = n3305_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4476_o = n3267_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4476_o = n3238_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4476_o = n3202_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4476_o = n3176_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4476_o = n3150_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4476_o = n3124_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4476_o = n3095_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4476_o = n3066_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4476_o = n3032_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4476_o = n3001_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4476_o = n2843_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4476_o = n2581_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4476_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4476_o = 1'b0;
      default: n4476_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4479_o = n2583_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4479_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4479_o = 1'b0;
      default: n4479_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4482_o = n4022_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4482_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4482_o = 1'b0;
      default: n4482_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4485_o = n2625_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4485_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4485_o = 1'b0;
      default: n4485_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4488_o = n2669_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4488_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4488_o = 1'b0;
      default: n4488_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4491_o = n4094_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4491_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4491_o = 1'b0;
      default: n4491_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4494_o = n4096_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4494_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4494_o = 1'b0;
      default: n4494_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4497_o = n2868_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4497_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4497_o = 1'b0;
      default: n4497_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4499_o = n3613_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4499_o = n3548_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4499_o = n3096_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4499_o = n2584_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4499_o = n2160_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4499_o = n2160_o;
      default: n4499_o = n2160_o;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4500_o = n3614_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4500_o = n3549_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4500_o = n3097_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4500_o = n2585_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4500_o = n2164_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4500_o = n2164_o;
      default: n4500_o = n2164_o;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4502_o = n3906_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4502_o = n3709_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4502_o = n2909_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4502_o = n2898_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4502_o = n2471_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4502_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4502_o = 1'b0;
      default: n4502_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4505_o = n4194_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4505_o = n3447_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4505_o = n3413_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4505_o = n2970_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4505_o = n2845_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4505_o = n2751_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4505_o = n2587_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4505_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4505_o = 1'b0;
      default: n4505_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4508_o = n3615_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4508_o = n3550_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4508_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4508_o = 1'b0;
      default: n4508_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4511_o = n3712_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4511_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4511_o = 1'b0;
      default: n4511_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4514_o = n3269_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4514_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4514_o = 1'b0;
      default: n4514_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4517_o = n2779_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4517_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4517_o = 1'b0;
      default: n4517_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4520_o = n2781_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4520_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4520_o = 1'b0;
      default: n4520_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4523_o = n2764_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4523_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4523_o = 1'b0;
      default: n4523_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4526_o = n2766_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4526_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4526_o = 1'b0;
      default: n4526_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4529_o = n4024_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4529_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4529_o = 1'b0;
      default: n4529_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4277_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4532_o = n2589_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4532_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4532_o = 1'b0;
      default: n4532_o = 1'b0;
    endcase
  /* decoder.vhd:2020:14  */
  assign n4536_o = ~res_i;
  /* decoder.vhd:2035:7  */
  assign n4539_o = bus_clear_f1_i ? 1'b0 : f1_q;
  /* decoder.vhd:2033:7  */
  assign n4541_o = bus_set_f1_i ? 1'b1 : n4539_o;
  /* decoder.vhd:2044:28  */
  assign n4543_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:2044:9  */
  assign n4545_o = n4543_o ? 1'b0 : branch_taken_q;
  /* decoder.vhd:2042:9  */
  assign n4547_o = branch_taken_s ? 1'b1 : n4545_o;
  /* decoder.vhd:2053:27  */
  assign n4548_o = ~f1_q;
  /* decoder.vhd:2052:9  */
  assign n4549_o = cpl_f1_s ? n4548_o : n4541_o;
  /* decoder.vhd:2050:9  */
  assign n4551_o = clear_f1_s ? 1'b0 : n4549_o;
  /* decoder.vhd:2059:9  */
  assign n4553_o = set_mb_s ? 1'b1 : mb_q;
  /* decoder.vhd:2057:9  */
  assign n4555_o = clear_mb_s ? 1'b0 : n4553_o;
  /* decoder.vhd:2039:7  */
  assign n4559_o = en_clk_i ? n4551_o : n4541_o;
  /* decoder.vhd:2039:7  */
  assign n4561_o = en_clk_i & ent0_clk_s;
  /* decoder.vhd:2115:27  */
  assign n4575_o = read_dec_s ? data_s : 8'b11111111;
  /* decoder.vhd:2117:48  */
  assign n4577_o = dm_write_dmem_s & en_clk_i;
  /* decoder.vhd:2118:48  */
  assign n4578_o = pm_inc_pc_s | add_inc_pc_s;
  /* decoder.vhd:2119:48  */
  assign n4579_o = pm_write_pmem_addr_s | add_write_pmem_addr_s;
  /* decoder.vhd:2121:48  */
  assign n4580_o = bus_read_bus_s | add_read_bus_s;
  /* decoder.vhd:305:5  */
  assign n4581_o = en_clk_i ? n1995_o : opc_opcode_q;
  /* decoder.vhd:305:5  */
  always @(posedge clk_i or posedge n1989_o)
    if (n1989_o)
      n4582_q <= 8'b00000000;
    else
      n4582_q <= n4581_o;
  /* decoder.vhd:2031:5  */
  assign n4583_o = en_clk_i ? n4547_o : branch_taken_q;
  /* decoder.vhd:2031:5  */
  always @(posedge clk_i or posedge n4536_o)
    if (n4536_o)
      n4584_q <= 1'b0;
    else
      n4584_q <= n4583_o;
  /* decoder.vhd:2031:5  */
  always @(posedge clk_i or posedge n4536_o)
    if (n4536_o)
      n4585_q <= 1'b0;
    else
      n4585_q <= n4559_o;
  /* decoder.vhd:2031:5  */
  assign n4586_o = en_clk_i ? n4555_o : mb_q;
  /* decoder.vhd:2031:5  */
  always @(posedge clk_i or posedge n4536_o)
    if (n4536_o)
      n4587_q <= 1'b0;
    else
      n4587_q <= n4586_o;
  /* decoder.vhd:2031:5  */
  assign n4588_o = n4561_o ? 1'b1 : t0_dir_q;
  /* decoder.vhd:2031:5  */
  always @(posedge clk_i or posedge n4536_o)
    if (n4536_o)
      n4589_q <= 1'b0;
    else
      n4589_q <= n4588_o;
  /* decoder.vhd:305:5  */
  assign n4590_o = en_clk_i ? n1996_o : mnemonic_q;
  /* decoder.vhd:305:5  */
  always @(posedge clk_i or posedge n1989_o)
    if (n1989_o)
      n4591_q <= 6'b101001;
    else
      n4591_q <= n4590_o;
  /* decoder.vhd:301:5  */
  assign n4592_o = {n4401_o, n4400_o};
endmodule

module upi41_db_bus_1
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_bus_i,
   input  read_bus_i,
   input  write_sts_i,
   input  f0_i,
   input  f1_i,
   input  ibf_int_i,
   input  en_dma_i,
   input  en_flags_i,
   input  write_p2_i,
   input  dack_n_i,
   input  a0_i,
   input  cs_n_i,
   input  rd_n_i,
   input  wr_n_i,
   input  [7:0] db_i,
   output [7:0] data_o,
   output set_f1_o,
   output clear_f1_o,
   output ibf_o,
   output obf_o,
   output int_n_o,
   output mint_ibf_n_o,
   output mint_obf_o,
   output dma_o,
   output drq_o,
   output [7:0] db_o,
   output db_dir_o);
  wire read_s;
  wire read_q;
  wire read_hold_q;
  wire write_s;
  wire write_q;
  wire read_pulse_s;
  wire write_pulse_s;
  wire a0_q;
  wire ibf_q;
  wire obf_q;
  wire [7:0] dbbin_q;
  wire [7:0] dbbout_q;
  wire [3:0] sts_q;
  wire dma_q;
  wire flags_q;
  wire ext_acc_s;
  wire dack_s;
  wire n1002_o;
  wire n1003_o;
  wire n1004_o;
  wire n1005_o;
  wire n1006_o;
  wire n1007_o;
  wire n1008_o;
  wire n1009_o;
  wire n1011_o;
  wire n1014_o;
  wire n1016_o;
  wire n1017_o;
  wire n1018_o;
  wire n1020_o;
  wire n1034_o;
  wire n1035_o;
  wire n1036_o;
  wire n1037_o;
  wire n1039_o;
  wire n1041_o;
  wire n1042_o;
  wire n1044_o;
  wire n1046_o;
  wire [7:0] n1047_o;
  wire n1048_o;
  wire n1049_o;
  wire n1051_o;
  wire [7:0] n1052_o;
  wire n1053_o;
  wire n1054_o;
  wire n1056_o;
  wire [3:0] n1057_o;
  wire [3:0] n1058_o;
  wire n1060_o;
  wire [3:0] n1061_o;
  wire n1062_o;
  wire n1064_o;
  wire [3:0] n1066_o;
  wire n1068_o;
  wire n1070_o;
  wire n1075_o;
  wire n1076_o;
  wire n1077_o;
  wire n1079_o;
  wire n1080_o;
  wire n1081_o;
  wire n1082_o;
  wire n1083_o;
  wire n1084_o;
  wire n1086_o;
  wire n1087_o;
  wire n1116_o;
  wire n1117_o;
  wire n1118_o;
  wire n1119_o;
  wire [7:0] n1120_o;
  wire [4:0] n1121_o;
  wire [5:0] n1122_o;
  wire [6:0] n1123_o;
  wire [7:0] n1124_o;
  wire [7:0] n1126_o;
  wire [4:0] n1128_o;
  wire [5:0] n1129_o;
  wire [6:0] n1130_o;
  wire [7:0] n1131_o;
  wire n1133_o;
  wire n1134_o;
  wire [7:0] n1136_o;
  wire n1139_o;
  wire n1140_o;
  wire n1143_o;
  wire n1144_o;
  wire n1145_o;
  reg n1147_q;
  reg n1148_q;
  reg n1149_q;
  reg n1150_q;
  reg n1151_q;
  reg n1152_q;
  reg [7:0] n1153_q;
  wire [7:0] n1154_o;
  reg [7:0] n1155_q;
  wire [3:0] n1156_o;
  reg [3:0] n1157_q;
  wire n1158_o;
  reg n1159_q;
  wire n1160_o;
  reg n1161_q;
  reg n1162_q;
  reg n1163_q;
  assign data_o = n1136_o;
  assign set_f1_o = n1116_o;
  assign clear_f1_o = n1118_o;
  assign ibf_o = ibf_q;
  assign obf_o = obf_q;
  assign int_n_o = n1162_q;
  assign mint_ibf_n_o = n1140_o;
  assign mint_obf_o = n1145_o;
  assign dma_o = dma_q;
  assign drq_o = n1163_q;
  assign db_o = n1120_o;
  assign db_dir_o = n1134_o;
  /* upi41_db_bus.vhd:103:10  */
  assign read_s = n1007_o; // (signal)
  /* upi41_db_bus.vhd:103:18  */
  assign read_q = n1147_q; // (signal)
  /* upi41_db_bus.vhd:104:10  */
  assign read_hold_q = n1148_q; // (signal)
  /* upi41_db_bus.vhd:105:10  */
  assign write_s = n1009_o; // (signal)
  /* upi41_db_bus.vhd:105:19  */
  assign write_q = n1149_q; // (signal)
  /* upi41_db_bus.vhd:106:10  */
  assign read_pulse_s = n1035_o; // (signal)
  /* upi41_db_bus.vhd:106:24  */
  assign write_pulse_s = n1037_o; // (signal)
  /* upi41_db_bus.vhd:108:10  */
  assign a0_q = n1150_q; // (signal)
  /* upi41_db_bus.vhd:110:10  */
  assign ibf_q = n1151_q; // (signal)
  /* upi41_db_bus.vhd:110:17  */
  assign obf_q = n1152_q; // (signal)
  /* upi41_db_bus.vhd:113:10  */
  assign dbbin_q = n1153_q; // (signal)
  /* upi41_db_bus.vhd:114:10  */
  assign dbbout_q = n1155_q; // (signal)
  /* upi41_db_bus.vhd:116:10  */
  assign sts_q = n1157_q; // (signal)
  /* upi41_db_bus.vhd:118:10  */
  assign dma_q = n1159_q; // (signal)
  /* upi41_db_bus.vhd:119:10  */
  assign flags_q = n1161_q; // (signal)
  /* upi41_db_bus.vhd:121:10  */
  assign ext_acc_s = n1005_o; // (signal)
  /* upi41_db_bus.vhd:122:10  */
  assign dack_s = n1003_o; // (signal)
  /* upi41_db_bus.vhd:142:25  */
  assign n1002_o = ~dack_n_i;
  /* upi41_db_bus.vhd:142:31  */
  assign n1003_o = n1002_o & dma_q;
  /* upi41_db_bus.vhd:143:23  */
  assign n1004_o = ~cs_n_i;
  /* upi41_db_bus.vhd:143:29  */
  assign n1005_o = n1004_o | dack_s;
  /* upi41_db_bus.vhd:144:37  */
  assign n1006_o = ~rd_n_i;
  /* upi41_db_bus.vhd:144:26  */
  assign n1007_o = ext_acc_s & n1006_o;
  /* upi41_db_bus.vhd:145:37  */
  assign n1008_o = ~wr_n_i;
  /* upi41_db_bus.vhd:145:26  */
  assign n1009_o = ext_acc_s & n1008_o;
  /* upi41_db_bus.vhd:149:14  */
  assign n1011_o = ~res_i;
  /* upi41_db_bus.vhd:161:7  */
  assign n1014_o = ext_acc_s ? 1'b0 : read_hold_q;
  /* upi41_db_bus.vhd:159:7  */
  assign n1016_o = read_s ? 1'b1 : n1014_o;
  /* upi41_db_bus.vhd:167:20  */
  assign n1017_o = read_s | write_s;
  /* upi41_db_bus.vhd:167:7  */
  assign n1018_o = n1017_o ? a0_i : a0_q;
  /* upi41_db_bus.vhd:165:7  */
  assign n1020_o = dack_s ? 1'b0 : n1018_o;
  /* upi41_db_bus.vhd:174:31  */
  assign n1034_o = ~read_s;
  /* upi41_db_bus.vhd:174:27  */
  assign n1035_o = read_q & n1034_o;
  /* upi41_db_bus.vhd:175:32  */
  assign n1036_o = ~write_s;
  /* upi41_db_bus.vhd:175:28  */
  assign n1037_o = write_q & n1036_o;
  /* upi41_db_bus.vhd:185:14  */
  assign n1039_o = ~res_i;
  /* upi41_db_bus.vhd:198:32  */
  assign n1041_o = ~a0_q;
  /* upi41_db_bus.vhd:198:23  */
  assign n1042_o = read_pulse_s & n1041_o;
  /* upi41_db_bus.vhd:200:7  */
  assign n1044_o = write_pulse_s ? 1'b0 : n1162_q;
  /* upi41_db_bus.vhd:200:7  */
  assign n1046_o = write_pulse_s ? 1'b1 : ibf_q;
  /* upi41_db_bus.vhd:200:7  */
  assign n1047_o = write_pulse_s ? db_i : dbbin_q;
  /* upi41_db_bus.vhd:198:7  */
  assign n1048_o = n1042_o ? n1162_q : n1044_o;
  /* upi41_db_bus.vhd:198:7  */
  assign n1049_o = n1042_o ? ibf_q : n1046_o;
  /* upi41_db_bus.vhd:198:7  */
  assign n1051_o = n1042_o ? 1'b0 : obf_q;
  /* upi41_db_bus.vhd:198:7  */
  assign n1052_o = n1042_o ? dbbin_q : n1047_o;
  /* upi41_db_bus.vhd:206:29  */
  assign n1053_o = read_s | write_s;
  /* upi41_db_bus.vhd:206:17  */
  assign n1054_o = dack_s & n1053_o;
  /* upi41_db_bus.vhd:206:7  */
  assign n1056_o = n1054_o ? 1'b0 : n1163_q;
  /* upi41_db_bus.vhd:217:29  */
  assign n1057_o = data_i[7:4];
  /* upi41_db_bus.vhd:216:9  */
  assign n1058_o = write_sts_i ? n1057_o : sts_q;
  /* upi41_db_bus.vhd:214:9  */
  assign n1060_o = read_bus_i ? 1'b0 : n1049_o;
  /* upi41_db_bus.vhd:214:9  */
  assign n1061_o = read_bus_i ? sts_q : n1058_o;
  /* upi41_db_bus.vhd:211:9  */
  assign n1062_o = write_bus_i ? n1049_o : n1060_o;
  /* upi41_db_bus.vhd:210:7  */
  assign n1064_o = n1083_o ? 1'b1 : n1051_o;
  /* upi41_db_bus.vhd:211:9  */
  assign n1066_o = write_bus_i ? sts_q : n1061_o;
  /* upi41_db_bus.vhd:210:7  */
  assign n1068_o = n1080_o ? 1'b1 : n1048_o;
  /* upi41_db_bus.vhd:225:11  */
  assign n1070_o = en_dma_i ? 1'b0 : n1056_o;
  /* upi41_db_bus.vhd:233:20  */
  assign n1075_o = dma_q & write_p2_i;
  /* upi41_db_bus.vhd:233:45  */
  assign n1076_o = data_i[6];
  /* upi41_db_bus.vhd:233:35  */
  assign n1077_o = n1075_o & n1076_o;
  /* upi41_db_bus.vhd:233:11  */
  assign n1079_o = n1077_o ? 1'b1 : n1070_o;
  /* upi41_db_bus.vhd:210:7  */
  assign n1080_o = en_clk_i & ibf_int_i;
  /* upi41_db_bus.vhd:210:7  */
  assign n1081_o = en_clk_i ? n1079_o : n1056_o;
  /* upi41_db_bus.vhd:210:7  */
  assign n1082_o = en_clk_i ? n1062_o : n1049_o;
  /* upi41_db_bus.vhd:210:7  */
  assign n1083_o = en_clk_i & write_bus_i;
  /* upi41_db_bus.vhd:210:7  */
  assign n1084_o = en_clk_i & write_bus_i;
  /* upi41_db_bus.vhd:210:7  */
  assign n1086_o = en_clk_i & en_dma_i;
  /* upi41_db_bus.vhd:210:7  */
  assign n1087_o = en_clk_i & en_flags_i;
  /* upi41_db_bus.vhd:250:31  */
  assign n1116_o = write_pulse_s & a0_q;
  /* upi41_db_bus.vhd:251:40  */
  assign n1117_o = ~a0_q;
  /* upi41_db_bus.vhd:251:31  */
  assign n1118_o = write_pulse_s & n1117_o;
  /* upi41_db_bus.vhd:254:36  */
  assign n1119_o = ~a0_q;
  /* upi41_db_bus.vhd:254:26  */
  assign n1120_o = n1119_o ? dbbout_q : n1126_o;
  /* upi41_db_bus.vhd:255:23  */
  assign n1121_o = {sts_q, f1_i};
  /* upi41_db_bus.vhd:255:30  */
  assign n1122_o = {n1121_o, f0_i};
  /* upi41_db_bus.vhd:255:37  */
  assign n1123_o = {n1122_o, ibf_q};
  /* upi41_db_bus.vhd:255:45  */
  assign n1124_o = {n1123_o, obf_q};
  /* upi41_db_bus.vhd:254:42  */
  assign n1126_o = 1'b1 ? n1124_o : n1131_o;
  /* upi41_db_bus.vhd:256:24  */
  assign n1128_o = {4'b0000, f1_i};
  /* upi41_db_bus.vhd:256:31  */
  assign n1129_o = {n1128_o, f0_i};
  /* upi41_db_bus.vhd:256:38  */
  assign n1130_o = {n1129_o, ibf_q};
  /* upi41_db_bus.vhd:256:46  */
  assign n1131_o = {n1130_o, obf_q};
  /* upi41_db_bus.vhd:257:36  */
  assign n1133_o = ext_acc_s & read_hold_q;
  /* upi41_db_bus.vhd:257:21  */
  assign n1134_o = n1133_o ? 1'b1 : 1'b0;
  /* upi41_db_bus.vhd:259:17  */
  assign n1136_o = read_bus_i ? dbbin_q : 8'b11111111;
  /* upi41_db_bus.vhd:262:36  */
  assign n1139_o = flags_q & ibf_q;
  /* upi41_db_bus.vhd:262:23  */
  assign n1140_o = n1139_o ? 1'b0 : 1'b1;
  /* upi41_db_bus.vhd:263:46  */
  assign n1143_o = ~obf_q;
  /* upi41_db_bus.vhd:263:36  */
  assign n1144_o = flags_q & n1143_o;
  /* upi41_db_bus.vhd:263:23  */
  assign n1145_o = n1144_o ? 1'b0 : 1'b1;
  /* upi41_db_bus.vhd:155:5  */
  always @(posedge clk_i or posedge n1011_o)
    if (n1011_o)
      n1147_q <= 1'b0;
    else
      n1147_q <= read_s;
  /* upi41_db_bus.vhd:155:5  */
  always @(posedge clk_i or posedge n1011_o)
    if (n1011_o)
      n1148_q <= 1'b0;
    else
      n1148_q <= n1016_o;
  /* upi41_db_bus.vhd:155:5  */
  always @(posedge clk_i or posedge n1011_o)
    if (n1011_o)
      n1149_q <= 1'b0;
    else
      n1149_q <= write_s;
  /* upi41_db_bus.vhd:155:5  */
  always @(posedge clk_i or posedge n1011_o)
    if (n1011_o)
      n1150_q <= 1'b0;
    else
      n1150_q <= n1020_o;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1151_q <= 1'b0;
    else
      n1151_q <= n1082_o;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1152_q <= 1'b0;
    else
      n1152_q <= n1064_o;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1153_q <= 8'b00000000;
    else
      n1153_q <= n1052_o;
  /* upi41_db_bus.vhd:196:5  */
  assign n1154_o = n1084_o ? data_i : dbbout_q;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1155_q <= 8'b00000000;
    else
      n1155_q <= n1154_o;
  /* upi41_db_bus.vhd:196:5  */
  assign n1156_o = en_clk_i ? n1066_o : sts_q;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1157_q <= 4'b0000;
    else
      n1157_q <= n1156_o;
  /* upi41_db_bus.vhd:196:5  */
  assign n1158_o = n1086_o ? 1'b1 : dma_q;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1159_q <= 1'b0;
    else
      n1159_q <= n1158_o;
  /* upi41_db_bus.vhd:196:5  */
  assign n1160_o = n1087_o ? 1'b1 : flags_q;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1161_q <= 1'b0;
    else
      n1161_q <= n1160_o;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1162_q <= 1'b1;
    else
      n1162_q <= n1068_o;
  /* upi41_db_bus.vhd:196:5  */
  always @(posedge clk_i or posedge n1039_o)
    if (n1039_o)
      n1163_q <= 1'b0;
    else
      n1163_q <= n1081_o;
endmodule

module t48_cond_branch
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  compute_take_i,
   input  [3:0] branch_cond_i,
   input  [7:0] accu_i,
   input  t0_i,
   input  t1_i,
   input  int_n_i,
   input  f0_i,
   input  f1_i,
   input  tf_i,
   input  carry_i,
   input  ibf_i,
   input  obf_i,
   input  [2:0] comp_value_i,
   output take_branch_o);
  wire take_branch_s;
  wire take_branch_q;
  wire n906_o;
  wire n908_o;
  wire n909_o;
  wire n911_o;
  wire n912_o;
  wire n913_o;
  wire n914_o;
  wire n915_o;
  wire n916_o;
  wire n917_o;
  wire n918_o;
  wire n919_o;
  wire n920_o;
  wire n921_o;
  wire n922_o;
  wire n923_o;
  wire n924_o;
  wire n925_o;
  wire n926_o;
  wire n927_o;
  wire n928_o;
  wire n930_o;
  wire n931_o;
  wire n932_o;
  wire n934_o;
  wire n936_o;
  wire n938_o;
  wire n939_o;
  wire n941_o;
  wire n942_o;
  wire n943_o;
  wire n945_o;
  wire n946_o;
  wire n947_o;
  wire n949_o;
  wire n951_o;
  wire n952_o;
  wire n954_o;
  wire n956_o;
  wire [10:0] n957_o;
  reg n959_o;
  wire n966_o;
  wire n969_o;
  wire n974_o;
  reg n975_q;
  wire n976_o;
  wire n977_o;
  wire n978_o;
  wire n979_o;
  wire n980_o;
  wire n981_o;
  wire n982_o;
  wire n983_o;
  wire [1:0] n984_o;
  reg n985_o;
  wire [1:0] n986_o;
  reg n987_o;
  wire n988_o;
  wire n989_o;
  assign take_branch_o = take_branch_q;
  /* cond_branch.vhd:90:10  */
  assign take_branch_s = n959_o; // (signal)
  /* cond_branch.vhd:91:10  */
  assign take_branch_q = n975_q; // (signal)
  /* cond_branch.vhd:119:9  */
  assign n906_o = n989_o ? 1'b1 : 1'b0;
  /* cond_branch.vhd:118:7  */
  assign n908_o = branch_cond_i == 4'b0000;
  /* cond_branch.vhd:126:33  */
  assign n909_o = accu_i[7];
  /* cond_branch.vhd:126:24  */
  assign n911_o = 1'b0 | n909_o;
  /* cond_branch.vhd:126:33  */
  assign n912_o = accu_i[6];
  /* cond_branch.vhd:126:24  */
  assign n913_o = n911_o | n912_o;
  /* cond_branch.vhd:126:33  */
  assign n914_o = accu_i[5];
  /* cond_branch.vhd:126:24  */
  assign n915_o = n913_o | n914_o;
  /* cond_branch.vhd:126:33  */
  assign n916_o = accu_i[4];
  /* cond_branch.vhd:126:24  */
  assign n917_o = n915_o | n916_o;
  /* cond_branch.vhd:126:33  */
  assign n918_o = accu_i[3];
  /* cond_branch.vhd:126:24  */
  assign n919_o = n917_o | n918_o;
  /* cond_branch.vhd:126:33  */
  assign n920_o = accu_i[2];
  /* cond_branch.vhd:126:24  */
  assign n921_o = n919_o | n920_o;
  /* cond_branch.vhd:126:33  */
  assign n922_o = accu_i[1];
  /* cond_branch.vhd:126:24  */
  assign n923_o = n921_o | n922_o;
  /* cond_branch.vhd:126:33  */
  assign n924_o = accu_i[0];
  /* cond_branch.vhd:126:24  */
  assign n925_o = n923_o | n924_o;
  /* cond_branch.vhd:128:49  */
  assign n926_o = comp_value_i[0];
  /* cond_branch.vhd:128:33  */
  assign n927_o = ~n926_o;
  /* cond_branch.vhd:128:31  */
  assign n928_o = n925_o == n927_o;
  /* cond_branch.vhd:124:7  */
  assign n930_o = branch_cond_i == 4'b0001;
  /* cond_branch.vhd:132:48  */
  assign n931_o = comp_value_i[0];
  /* cond_branch.vhd:132:34  */
  assign n932_o = carry_i == n931_o;
  /* cond_branch.vhd:131:7  */
  assign n934_o = branch_cond_i == 4'b0010;
  /* cond_branch.vhd:135:7  */
  assign n936_o = branch_cond_i == 4'b0011;
  /* cond_branch.vhd:139:7  */
  assign n938_o = branch_cond_i == 4'b0100;
  /* cond_branch.vhd:144:34  */
  assign n939_o = ~int_n_i;
  /* cond_branch.vhd:143:7  */
  assign n941_o = branch_cond_i == 4'b0101;
  /* cond_branch.vhd:148:45  */
  assign n942_o = comp_value_i[0];
  /* cond_branch.vhd:148:31  */
  assign n943_o = t0_i == n942_o;
  /* cond_branch.vhd:147:7  */
  assign n945_o = branch_cond_i == 4'b0110;
  /* cond_branch.vhd:152:45  */
  assign n946_o = comp_value_i[0];
  /* cond_branch.vhd:152:31  */
  assign n947_o = t1_i == n946_o;
  /* cond_branch.vhd:151:7  */
  assign n949_o = branch_cond_i == 4'b0111;
  /* cond_branch.vhd:155:7  */
  assign n951_o = branch_cond_i == 4'b1000;
  /* cond_branch.vhd:160:32  */
  assign n952_o = ~ibf_i;
  /* cond_branch.vhd:159:7  */
  assign n954_o = branch_cond_i == 4'b1001;
  /* cond_branch.vhd:163:7  */
  assign n956_o = branch_cond_i == 4'b1010;
  /* clock_ctrl.vhd:206:5  */
  assign n957_o = {n956_o, n954_o, n951_o, n949_o, n945_o, n941_o, n938_o, n936_o, n934_o, n930_o, n908_o};
  /* cond_branch.vhd:116:5  */
  always @*
    case (n957_o)
      11'b10000000000: n959_o = obf_i;
      11'b01000000000: n959_o = n952_o;
      11'b00100000000: n959_o = tf_i;
      11'b00010000000: n959_o = n947_o;
      11'b00001000000: n959_o = n943_o;
      11'b00000100000: n959_o = n939_o;
      11'b00000010000: n959_o = f1_i;
      11'b00000001000: n959_o = f0_i;
      11'b00000000100: n959_o = n932_o;
      11'b00000000010: n959_o = n928_o;
      11'b00000000001: n959_o = n906_o;
      default: n959_o = 1'b0;
    endcase
  /* cond_branch.vhd:188:14  */
  assign n966_o = ~res_i;
  /* cond_branch.vhd:192:7  */
  assign n969_o = en_clk_i & compute_take_i;
  /* cond_branch.vhd:191:5  */
  assign n974_o = n969_o ? take_branch_s : take_branch_q;
  /* cond_branch.vhd:191:5  */
  always @(posedge clk_i or posedge n966_o)
    if (n966_o)
      n975_q <= 1'b0;
    else
      n975_q <= n974_o;
  /* cond_branch.vhd:64:5  */
  assign n976_o = accu_i[0];
  assign n977_o = accu_i[1];
  /* cond_branch.vhd:191:5  */
  assign n978_o = accu_i[2];
  /* cond_branch.vhd:186:3  */
  assign n979_o = accu_i[3];
  assign n980_o = accu_i[4];
  assign n981_o = accu_i[5];
  /* cond_branch.vhd:116:5  */
  assign n982_o = accu_i[6];
  assign n983_o = accu_i[7];
  /* cond_branch.vhd:119:18  */
  assign n984_o = comp_value_i[1:0];
  /* cond_branch.vhd:119:18  */
  always @*
    case (n984_o)
      2'b00: n985_o = n976_o;
      2'b01: n985_o = n977_o;
      2'b10: n985_o = n978_o;
      2'b11: n985_o = n979_o;
    endcase
  /* cond_branch.vhd:119:18  */
  assign n986_o = comp_value_i[1:0];
  /* cond_branch.vhd:119:18  */
  always @*
    case (n986_o)
      2'b00: n987_o = n980_o;
      2'b01: n987_o = n981_o;
      2'b10: n987_o = n982_o;
      2'b11: n987_o = n983_o;
    endcase
  /* cond_branch.vhd:119:18  */
  assign n988_o = comp_value_i[2];
  /* cond_branch.vhd:119:18  */
  assign n989_o = n988_o ? n987_o : n985_o;
endmodule

module t48_clock_ctrl_1
  (input  clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  res_i,
   input  en_clk_i,
   input  multi_cycle_i,
   input  assert_psen_i,
   input  assert_prog_i,
   input  assert_rd_i,
   input  assert_wr_i,
   output xtal3_o,
   output t0_o,
   output [2:0] mstate_o,
   output second_cycle_o,
   output ale_o,
   output psen_o,
   output prog_o,
   output rd_o,
   output wr_o);
  wire [1:0] xtal_q;
  wire xtal2_s;
  wire xtal3_s;
  wire x2_s;
  wire x3_s;
  wire t0_q;
  wire [2:0] mstate_q;
  wire ale_q;
  wire psen_q;
  wire prog_q;
  wire rd_q;
  wire wr_q;
  wire second_cycle_q;
  wire multi_cycle_q;
  wire n682_o;
  wire n685_o;
  wire [1:0] n687_o;
  wire [1:0] n689_o;
  wire n692_o;
  wire n710_o;
  wire n711_o;
  wire n712_o;
  wire n716_o;
  wire n717_o;
  wire n718_o;
  wire n735_o;
  wire n743_o;
  wire n745_o;
  wire n747_o;
  wire n748_o;
  wire n750_o;
  wire n752_o;
  wire n753_o;
  wire n754_o;
  wire n756_o;
  wire n758_o;
  wire n760_o;
  wire n762_o;
  wire n764_o;
  wire n766_o;
  wire n768_o;
  wire n770_o;
  wire n772_o;
  wire n774_o;
  wire n775_o;
  wire n776_o;
  wire n777_o;
  wire n778_o;
  wire n779_o;
  wire n781_o;
  wire n783_o;
  wire n785_o;
  wire [4:0] n786_o;
  reg n788_o;
  reg n790_o;
  reg n792_o;
  reg n794_o;
  reg n796_o;
  wire n814_o;
  wire n817_o;
  wire n819_o;
  wire n821_o;
  wire n823_o;
  wire n825_o;
  wire [4:0] n826_o;
  reg [2:0] n833_o;
  wire n842_o;
  wire n845_o;
  wire n847_o;
  wire n848_o;
  wire n850_o;
  wire n851_o;
  wire n853_o;
  wire n854_o;
  wire n855_o;
  wire n857_o;
  wire n859_o;
  wire [1:0] n883_o;
  reg [1:0] n884_q;
  wire n885_o;
  reg n886_q;
  wire [2:0] n887_o;
  reg [2:0] n888_q;
  reg n889_q;
  reg n890_q;
  reg n891_q;
  reg n892_q;
  reg n893_q;
  wire n894_o;
  reg n895_q;
  wire n896_o;
  reg n897_q;
  assign xtal3_o = xtal3_s;
  assign t0_o = t0_q;
  assign mstate_o = mstate_q;
  assign second_cycle_o = second_cycle_q;
  assign ale_o = ale_q;
  assign psen_o = psen_q;
  assign prog_o = prog_q;
  assign rd_o = rd_q;
  assign wr_o = wr_q;
  /* clock_ctrl.vhd:90:10  */
  assign xtal_q = n884_q; // (signal)
  /* clock_ctrl.vhd:92:10  */
  assign xtal2_s = n735_o; // (signal)
  /* clock_ctrl.vhd:93:10  */
  assign xtal3_s = n743_o; // (signal)
  /* clock_ctrl.vhd:95:10  */
  assign x2_s = n712_o; // (signal)
  /* clock_ctrl.vhd:96:10  */
  assign x3_s = n718_o; // (signal)
  /* clock_ctrl.vhd:98:10  */
  assign t0_q = n886_q; // (signal)
  /* clock_ctrl.vhd:102:10  */
  assign mstate_q = n888_q; // (signal)
  /* clock_ctrl.vhd:104:10  */
  assign ale_q = n889_q; // (signal)
  /* clock_ctrl.vhd:105:10  */
  assign psen_q = n890_q; // (signal)
  /* clock_ctrl.vhd:106:10  */
  assign prog_q = n891_q; // (signal)
  /* clock_ctrl.vhd:107:10  */
  assign rd_q = n892_q; // (signal)
  /* clock_ctrl.vhd:108:10  */
  assign wr_q = n893_q; // (signal)
  /* clock_ctrl.vhd:112:10  */
  assign second_cycle_q = n895_q; // (signal)
  /* clock_ctrl.vhd:113:10  */
  assign multi_cycle_q = n897_q; // (signal)
  /* clock_ctrl.vhd:137:16  */
  assign n682_o = ~res_i;
  /* clock_ctrl.vhd:143:21  */
  assign n685_o = $unsigned(xtal_q) < $unsigned(2'b10);
  /* clock_ctrl.vhd:144:30  */
  assign n687_o = xtal_q + 2'b01;
  /* clock_ctrl.vhd:143:11  */
  assign n689_o = n685_o ? n687_o : 2'b00;
  /* clock_ctrl.vhd:149:11  */
  assign n692_o = xtal3_s ? 1'b1 : 1'b0;
  /* clock_ctrl.vhd:164:25  */
  assign n710_o = xtal_q == 2'b01;
  /* clock_ctrl.vhd:164:29  */
  assign n711_o = n710_o & xtal_en_i;
  /* clock_ctrl.vhd:164:13  */
  assign n712_o = n711_o ? 1'b1 : 1'b0;
  /* clock_ctrl.vhd:167:25  */
  assign n716_o = xtal_q == 2'b10;
  /* clock_ctrl.vhd:167:29  */
  assign n717_o = n716_o & xtal_en_i;
  /* clock_ctrl.vhd:167:13  */
  assign n718_o = n717_o ? 1'b1 : 1'b0;
  /* t48_pack-p.vhd:75:5  */
  assign n735_o = x2_s ? 1'b1 : 1'b0;
  /* t48_pack-p.vhd:75:5  */
  assign n743_o = x3_s ? 1'b1 : 1'b0;
  /* clock_ctrl.vhd:206:14  */
  assign n745_o = ~res_i;
  /* clock_ctrl.vhd:218:26  */
  assign n747_o = ~second_cycle_q;
  /* clock_ctrl.vhd:218:22  */
  assign n748_o = xtal2_s & n747_o;
  /* clock_ctrl.vhd:218:11  */
  assign n750_o = n753_o ? 1'b1 : rd_q;
  /* clock_ctrl.vhd:218:11  */
  assign n752_o = n754_o ? 1'b1 : wr_q;
  /* clock_ctrl.vhd:218:11  */
  assign n753_o = n748_o & assert_rd_i;
  /* clock_ctrl.vhd:218:11  */
  assign n754_o = n748_o & assert_wr_i;
  /* clock_ctrl.vhd:216:9  */
  assign n756_o = mstate_q == 3'b100;
  /* clock_ctrl.vhd:228:11  */
  assign n758_o = xtal3_s ? 1'b0 : psen_q;
  /* clock_ctrl.vhd:227:9  */
  assign n760_o = mstate_q == 3'b000;
  /* clock_ctrl.vhd:233:11  */
  assign n762_o = xtal3_s ? 1'b0 : prog_q;
  /* clock_ctrl.vhd:233:11  */
  assign n764_o = xtal3_s ? 1'b0 : rd_q;
  /* clock_ctrl.vhd:233:11  */
  assign n766_o = xtal3_s ? 1'b0 : wr_q;
  /* clock_ctrl.vhd:232:9  */
  assign n768_o = mstate_q == 3'b001;
  /* clock_ctrl.vhd:243:11  */
  assign n770_o = xtal3_s ? 1'b1 : ale_q;
  /* clock_ctrl.vhd:241:9  */
  assign n772_o = mstate_q == 3'b010;
  /* clock_ctrl.vhd:248:11  */
  assign n774_o = n775_o ? 1'b1 : psen_q;
  /* clock_ctrl.vhd:248:11  */
  assign n775_o = xtal3_s & assert_psen_i;
  /* clock_ctrl.vhd:257:22  */
  assign n776_o = xtal3_s & multi_cycle_q;
  /* clock_ctrl.vhd:258:32  */
  assign n777_o = ~second_cycle_q;
  /* clock_ctrl.vhd:258:28  */
  assign n778_o = n776_o & n777_o;
  /* clock_ctrl.vhd:258:51  */
  assign n779_o = n778_o & assert_prog_i;
  /* clock_ctrl.vhd:257:11  */
  assign n781_o = n779_o ? 1'b1 : prog_q;
  /* clock_ctrl.vhd:263:11  */
  assign n783_o = xtal2_s ? 1'b0 : ale_q;
  /* clock_ctrl.vhd:247:9  */
  assign n785_o = mstate_q == 3'b011;
  assign n786_o = {n785_o, n772_o, n768_o, n760_o, n756_o};
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n786_o)
      5'b10000: n788_o = n783_o;
      5'b01000: n788_o = n770_o;
      5'b00100: n788_o = ale_q;
      5'b00010: n788_o = ale_q;
      5'b00001: n788_o = ale_q;
      default: n788_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n786_o)
      5'b10000: n790_o = n774_o;
      5'b01000: n790_o = psen_q;
      5'b00100: n790_o = psen_q;
      5'b00010: n790_o = n758_o;
      5'b00001: n790_o = psen_q;
      default: n790_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n786_o)
      5'b10000: n792_o = n781_o;
      5'b01000: n792_o = prog_q;
      5'b00100: n792_o = n762_o;
      5'b00010: n792_o = prog_q;
      5'b00001: n792_o = prog_q;
      default: n792_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n786_o)
      5'b10000: n794_o = rd_q;
      5'b01000: n794_o = rd_q;
      5'b00100: n794_o = n764_o;
      5'b00010: n794_o = rd_q;
      5'b00001: n794_o = n750_o;
      default: n794_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n786_o)
      5'b10000: n796_o = wr_q;
      5'b01000: n796_o = wr_q;
      5'b00100: n796_o = n766_o;
      5'b00010: n796_o = wr_q;
      5'b00001: n796_o = n752_o;
      default: n796_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:292:14  */
  assign n814_o = ~res_i;
  /* clock_ctrl.vhd:303:11  */
  assign n817_o = mstate_q == 3'b100;
  /* clock_ctrl.vhd:306:11  */
  assign n819_o = mstate_q == 3'b000;
  /* clock_ctrl.vhd:309:11  */
  assign n821_o = mstate_q == 3'b001;
  /* clock_ctrl.vhd:312:11  */
  assign n823_o = mstate_q == 3'b010;
  /* clock_ctrl.vhd:315:11  */
  assign n825_o = mstate_q == 3'b011;
  assign n826_o = {n825_o, n823_o, n821_o, n819_o, n817_o};
  /* clock_ctrl.vhd:302:9  */
  always @*
    case (n826_o)
      5'b10000: n833_o = 3'b100;
      5'b01000: n833_o = 3'b011;
      5'b00100: n833_o = 3'b010;
      5'b00010: n833_o = 3'b001;
      5'b00001: n833_o = 3'b000;
      default: n833_o = 3'b000;
    endcase
  /* clock_ctrl.vhd:349:14  */
  assign n842_o = ~res_i;
  /* clock_ctrl.vhd:356:30  */
  assign n845_o = mstate_q == 3'b001;
  /* clock_ctrl.vhd:357:30  */
  assign n847_o = mstate_q == 3'b100;
  /* clock_ctrl.vhd:360:21  */
  assign n848_o = n845_o & multi_cycle_i;
  /* clock_ctrl.vhd:360:9  */
  assign n850_o = n848_o ? 1'b1 : multi_cycle_q;
  /* clock_ctrl.vhd:365:26  */
  assign n851_o = multi_cycle_q & n847_o;
  /* clock_ctrl.vhd:365:9  */
  assign n853_o = n851_o ? 1'b1 : second_cycle_q;
  /* clock_ctrl.vhd:371:27  */
  assign n854_o = multi_cycle_q & second_cycle_q;
  /* clock_ctrl.vhd:370:21  */
  assign n855_o = n847_o & n854_o;
  /* clock_ctrl.vhd:370:9  */
  assign n857_o = n855_o ? 1'b0 : n853_o;
  /* clock_ctrl.vhd:370:9  */
  assign n859_o = n855_o ? 1'b0 : n850_o;
  /* clock_ctrl.vhd:141:7  */
  assign n883_o = xtal_en_i ? n689_o : xtal_q;
  /* clock_ctrl.vhd:141:7  */
  always @(posedge xtal_i or posedge n682_o)
    if (n682_o)
      n884_q <= 2'b00;
    else
      n884_q <= n883_o;
  /* clock_ctrl.vhd:141:7  */
  assign n885_o = xtal_en_i ? n692_o : t0_q;
  /* clock_ctrl.vhd:141:7  */
  always @(posedge xtal_i or posedge n682_o)
    if (n682_o)
      n886_q <= 1'b0;
    else
      n886_q <= n885_o;
  /* clock_ctrl.vhd:299:5  */
  assign n887_o = en_clk_i ? n833_o : mstate_q;
  /* clock_ctrl.vhd:299:5  */
  always @(posedge clk_i or posedge n814_o)
    if (n814_o)
      n888_q <= 3'b010;
    else
      n888_q <= n887_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n745_o)
    if (n745_o)
      n889_q <= 1'b0;
    else
      n889_q <= n788_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n745_o)
    if (n745_o)
      n890_q <= 1'b0;
    else
      n890_q <= n790_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n745_o)
    if (n745_o)
      n891_q <= 1'b0;
    else
      n891_q <= n792_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n745_o)
    if (n745_o)
      n892_q <= 1'b0;
    else
      n892_q <= n794_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n745_o)
    if (n745_o)
      n893_q <= 1'b0;
    else
      n893_q <= n796_o;
  /* clock_ctrl.vhd:353:5  */
  assign n894_o = en_clk_i ? n857_o : second_cycle_q;
  /* clock_ctrl.vhd:353:5  */
  always @(posedge clk_i or posedge n842_o)
    if (n842_o)
      n895_q <= 1'b0;
    else
      n895_q <= n894_o;
  /* clock_ctrl.vhd:353:5  */
  assign n896_o = en_clk_i ? n859_o : multi_cycle_q;
  /* clock_ctrl.vhd:353:5  */
  always @(posedge clk_i or posedge n842_o)
    if (n842_o)
      n897_q <= 1'b0;
    else
      n897_q <= n896_o;
endmodule

module t48_bus_mux
  (input  [7:0] alu_data_i,
   input  [7:0] bus_data_i,
   input  [7:0] dec_data_i,
   input  [7:0] dm_data_i,
   input  [7:0] pm_data_i,
   input  [7:0] p1_data_i,
   input  [7:0] p2_data_i,
   input  [7:0] psw_data_i,
   input  [7:0] tim_data_i,
   output [7:0] data_o);
  wire [7:0] n664_o;
  wire [7:0] n665_o;
  wire [7:0] n666_o;
  wire [7:0] n667_o;
  wire [7:0] n668_o;
  wire [7:0] n669_o;
  wire [7:0] n670_o;
  wire [7:0] n671_o;
  assign data_o = n671_o;
  /* bus_mux.vhd:89:26  */
  assign n664_o = alu_data_i & bus_data_i;
  /* bus_mux.vhd:90:26  */
  assign n665_o = n664_o & dec_data_i;
  /* bus_mux.vhd:91:26  */
  assign n666_o = n665_o & dm_data_i;
  /* bus_mux.vhd:92:26  */
  assign n667_o = n666_o & pm_data_i;
  /* bus_mux.vhd:93:26  */
  assign n668_o = n667_o & p1_data_i;
  /* bus_mux.vhd:94:26  */
  assign n669_o = n668_o & p2_data_i;
  /* bus_mux.vhd:95:26  */
  assign n670_o = n669_o & psw_data_i;
  /* bus_mux.vhd:96:26  */
  assign n671_o = n670_o & tim_data_i;
endmodule

module t48_alu
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_accu_i,
   input  write_shadow_i,
   input  write_temp_reg_i,
   input  read_alu_i,
   input  carry_i,
   input  [3:0] alu_op_i,
   input  use_carry_i,
   input  da_high_i,
   input  accu_low_i,
   input  p06_temp_reg_i,
   input  p60_temp_reg_i,
   output [7:0] data_o,
   output carry_o,
   output aux_carry_o,
   output da_overflow_o);
  wire [7:0] accumulator_q;
  wire [7:0] accu_shadow_q;
  wire [7:0] temp_req_q;
  wire [7:0] in_a_s;
  wire [7:0] in_b_s;
  wire [7:0] data_s;
  wire [8:0] add_result_s;
  wire n413_o;
  wire [3:0] n415_o;
  wire [3:0] n416_o;
  wire [3:0] n417_o;
  wire [3:0] n418_o;
  wire [3:0] n419_o;
  wire [3:0] n420_o;
  wire [7:0] n421_o;
  wire [7:0] n423_o;
  wire [7:0] n424_o;
  wire [7:0] n426_o;
  wire [7:0] n428_o;
  wire n429_o;
  wire [7:0] n443_o;
  wire n445_o;
  wire [7:0] n446_o;
  wire n448_o;
  wire [7:0] n449_o;
  wire n451_o;
  wire [7:0] n452_o;
  wire n453_o;
  wire n455_o;
  wire [7:0] n456_o;
  wire n458_o;
  wire n460_o;
  wire [6:0] n461_o;
  wire n462_o;
  wire n463_o;
  wire n464_o;
  wire n466_o;
  wire [6:0] n467_o;
  wire n468_o;
  wire n469_o;
  wire n470_o;
  wire n472_o;
  wire [3:0] n473_o;
  wire [3:0] n474_o;
  wire n476_o;
  wire [7:0] n477_o;
  wire n479_o;
  wire [7:0] n480_o;
  wire n482_o;
  wire [3:0] n483_o;
  wire [3:0] n484_o;
  wire [7:0] n485_o;
  wire n487_o;
  wire n489_o;
  wire [12:0] n490_o;
  reg n492_o;
  wire n494_o;
  wire n495_o;
  wire n496_o;
  wire n497_o;
  wire n498_o;
  wire n500_o;
  wire n501_o;
  wire n502_o;
  wire n503_o;
  wire n504_o;
  wire n505_o;
  reg n507_o;
  wire [2:0] n508_o;
  wire [2:0] n509_o;
  wire [2:0] n510_o;
  wire [2:0] n511_o;
  wire [2:0] n512_o;
  wire [2:0] n514_o;
  wire [2:0] n515_o;
  wire [2:0] n516_o;
  wire [2:0] n517_o;
  wire [2:0] n518_o;
  wire [2:0] n519_o;
  wire [2:0] n520_o;
  reg [2:0] n522_o;
  wire [2:0] n523_o;
  wire [2:0] n524_o;
  wire [2:0] n525_o;
  wire [2:0] n526_o;
  wire [2:0] n527_o;
  wire [2:0] n529_o;
  wire [2:0] n530_o;
  wire [2:0] n531_o;
  wire [2:0] n532_o;
  wire [2:0] n533_o;
  wire [2:0] n534_o;
  wire [2:0] n535_o;
  reg [2:0] n537_o;
  wire n538_o;
  wire n539_o;
  wire n540_o;
  wire n541_o;
  wire n542_o;
  wire n544_o;
  wire n545_o;
  wire n546_o;
  wire n547_o;
  wire n548_o;
  wire n549_o;
  reg n551_o;
  wire n563_o;
  wire n566_o;
  localparam [8:0] n567_o = 9'b000000000;
  wire [7:0] n568_o;
  wire [8:0] n570_o;
  wire [8:0] n572_o;
  localparam [8:0] n574_o = 9'b000000000;
  wire [7:0] n575_o;
  wire n577_o;
  wire n579_o;
  wire [1:0] n580_o;
  wire n582_o;
  reg n583_o;
  wire [7:0] n585_o;
  reg [7:0] n586_o;
  wire [8:0] n588_o;
  wire [8:0] n589_o;
  wire [8:0] n590_o;
  wire [8:0] n591_o;
  wire n592_o;
  wire n593_o;
  wire [1:0] n594_o;
  wire n595_o;
  wire n598_o;
  wire n600_o;
  wire n602_o;
  wire n603_o;
  wire n604_o;
  wire n605_o;
  wire n608_o;
  wire n610_o;
  wire n612_o;
  wire n613_o;
  wire [1:0] n614_o;
  reg n616_o;
  wire [3:0] n623_o;
  wire [3:0] n624_o;
  wire [3:0] n625_o;
  wire n633_o;
  wire n635_o;
  wire n636_o;
  wire n638_o;
  wire n639_o;
  wire n641_o;
  wire n642_o;
  wire n644_o;
  wire n645_o;
  wire n647_o;
  wire n648_o;
  reg n651_o;
  wire [7:0] n654_o;
  wire [7:0] n656_o;
  reg [7:0] n657_q;
  wire [7:0] n658_o;
  reg [7:0] n659_q;
  wire [7:0] n660_o;
  reg [7:0] n661_q;
  wire [7:0] n662_o;
  assign data_o = n654_o;
  assign carry_o = n492_o;
  assign aux_carry_o = n616_o;
  assign da_overflow_o = n651_o;
  /* alu.vhd:99:10  */
  assign accumulator_q = n657_q; // (signal)
  /* alu.vhd:100:10  */
  assign accu_shadow_q = n659_q; // (signal)
  /* alu.vhd:101:10  */
  assign temp_req_q = n661_q; // (signal)
  /* alu.vhd:103:10  */
  assign in_a_s = accu_shadow_q; // (signal)
  /* alu.vhd:104:10  */
  assign in_b_s = temp_req_q; // (signal)
  /* alu.vhd:106:10  */
  assign data_s = n662_o; // (signal)
  /* alu.vhd:108:10  */
  assign add_result_s = n591_o; // (signal)
  /* alu.vhd:122:14  */
  assign n413_o = ~res_i;
  /* alu.vhd:132:52  */
  assign n415_o = data_i[3:0];
  /* upi41_core.vhd:562:24  */
  assign n416_o = data_i[3:0];
  /* alu.vhd:131:11  */
  assign n417_o = accu_low_i ? n415_o : n416_o;
  /* upi41_core.vhd:545:3  */
  assign n418_o = data_i[7:4];
  /* upi41_core.vhd:545:3  */
  assign n419_o = accumulator_q[7:4];
  /* alu.vhd:131:11  */
  assign n420_o = accu_low_i ? n419_o : n418_o;
  /* upi41_core.vhd:545:3  */
  assign n421_o = {n420_o, n417_o};
  /* alu.vhd:138:9  */
  assign n423_o = write_shadow_i ? data_i : accumulator_q;
  /* alu.vhd:152:9  */
  assign n424_o = write_temp_reg_i ? data_i : temp_req_q;
  /* alu.vhd:149:9  */
  assign n426_o = p60_temp_reg_i ? 8'b01100000 : n424_o;
  /* alu.vhd:146:9  */
  assign n428_o = p06_temp_reg_i ? 8'b00000110 : n426_o;
  /* alu.vhd:128:7  */
  assign n429_o = en_clk_i & write_accu_i;
  /* alu.vhd:203:26  */
  assign n443_o = in_a_s & in_b_s;
  /* alu.vhd:202:7  */
  assign n445_o = alu_op_i == 4'b0000;
  /* alu.vhd:207:26  */
  assign n446_o = in_a_s | in_b_s;
  /* alu.vhd:206:7  */
  assign n448_o = alu_op_i == 4'b0001;
  /* alu.vhd:211:26  */
  assign n449_o = in_a_s ^ in_b_s;
  /* alu.vhd:210:7  */
  assign n451_o = alu_op_i == 4'b0010;
  /* alu.vhd:215:32  */
  assign n452_o = add_result_s[7:0];
  /* alu.vhd:216:32  */
  assign n453_o = add_result_s[8];
  /* alu.vhd:214:7  */
  assign n455_o = alu_op_i == 4'b1010;
  /* alu.vhd:220:19  */
  assign n456_o = ~in_a_s;
  /* alu.vhd:219:7  */
  assign n458_o = alu_op_i == 4'b0011;
  /* alu.vhd:223:7  */
  assign n460_o = alu_op_i == 4'b0100;
  /* alu.vhd:228:37  */
  assign n461_o = in_a_s[6:0];
  /* alu.vhd:229:37  */
  assign n462_o = in_a_s[7];
  /* alu.vhd:234:37  */
  assign n463_o = in_a_s[7];
  /* alu.vhd:231:9  */
  assign n464_o = use_carry_i ? carry_i : n463_o;
  /* alu.vhd:227:7  */
  assign n466_o = alu_op_i == 4'b0101;
  /* alu.vhd:239:37  */
  assign n467_o = in_a_s[7:1];
  /* alu.vhd:240:37  */
  assign n468_o = in_a_s[0];
  /* alu.vhd:245:37  */
  assign n469_o = in_a_s[0];
  /* alu.vhd:242:9  */
  assign n470_o = use_carry_i ? carry_i : n469_o;
  /* alu.vhd:238:7  */
  assign n472_o = alu_op_i == 4'b0110;
  /* alu.vhd:250:37  */
  assign n473_o = in_a_s[7:4];
  /* alu.vhd:251:37  */
  assign n474_o = in_a_s[3:0];
  /* alu.vhd:249:7  */
  assign n476_o = alu_op_i == 4'b0111;
  /* alu.vhd:255:31  */
  assign n477_o = add_result_s[7:0];
  /* alu.vhd:254:7  */
  assign n479_o = alu_op_i == 4'b1000;
  /* alu.vhd:259:31  */
  assign n480_o = add_result_s[7:0];
  /* alu.vhd:258:7  */
  assign n482_o = alu_op_i == 4'b1001;
  /* alu.vhd:263:25  */
  assign n483_o = in_b_s[7:4];
  /* alu.vhd:263:46  */
  assign n484_o = in_a_s[3:0];
  /* alu.vhd:263:38  */
  assign n485_o = {n483_o, n484_o};
  /* alu.vhd:262:7  */
  assign n487_o = alu_op_i == 4'b1011;
  /* alu.vhd:266:7  */
  assign n489_o = alu_op_i == 4'b1100;
  /* upi41_core.vhd:426:33  */
  assign n490_o = {n489_o, n487_o, n482_o, n479_o, n476_o, n472_o, n466_o, n460_o, n458_o, n455_o, n451_o, n448_o, n445_o};
  /* alu.vhd:200:5  */
  always @*
    case (n490_o)
      13'b1000000000000: n492_o = 1'b0;
      13'b0100000000000: n492_o = 1'b0;
      13'b0010000000000: n492_o = 1'b0;
      13'b0001000000000: n492_o = 1'b0;
      13'b0000100000000: n492_o = 1'b0;
      13'b0000010000000: n492_o = n468_o;
      13'b0000001000000: n492_o = n462_o;
      13'b0000000100000: n492_o = 1'b0;
      13'b0000000010000: n492_o = 1'b0;
      13'b0000000001000: n492_o = n453_o;
      13'b0000000000100: n492_o = 1'b0;
      13'b0000000000010: n492_o = 1'b0;
      13'b0000000000001: n492_o = 1'b0;
      default: n492_o = 1'b0;
    endcase
  /* upi41_core.vhd:422:33  */
  assign n494_o = n443_o[0];
  /* upi41_core.vhd:421:33  */
  assign n495_o = n446_o[0];
  /* upi41_core.vhd:420:33  */
  assign n496_o = n449_o[0];
  /* upi41_core.vhd:417:33  */
  assign n497_o = n452_o[0];
  /* upi41_core.vhd:416:33  */
  assign n498_o = n456_o[0];
  /* upi41_core.vhd:414:33  */
  assign n500_o = n467_o[0];
  /* upi41_core.vhd:413:33  */
  assign n501_o = n473_o[0];
  /* upi41_core.vhd:412:33  */
  assign n502_o = n477_o[0];
  /* upi41_core.vhd:411:33  */
  assign n503_o = n480_o[0];
  /* upi41_core.vhd:394:3  */
  assign n504_o = n485_o[0];
  /* upi41_core.vhd:394:3  */
  assign n505_o = in_a_s[0];
  /* alu.vhd:200:5  */
  always @*
    case (n490_o)
      13'b1000000000000: n507_o = n505_o;
      13'b0100000000000: n507_o = n504_o;
      13'b0010000000000: n507_o = n503_o;
      13'b0001000000000: n507_o = n502_o;
      13'b0000100000000: n507_o = n501_o;
      13'b0000010000000: n507_o = n500_o;
      13'b0000001000000: n507_o = n464_o;
      13'b0000000100000: n507_o = 1'b0;
      13'b0000000010000: n507_o = n498_o;
      13'b0000000001000: n507_o = n497_o;
      13'b0000000000100: n507_o = n496_o;
      13'b0000000000010: n507_o = n495_o;
      13'b0000000000001: n507_o = n494_o;
      default: n507_o = 1'b0;
    endcase
  /* upi41_core.vhd:394:3  */
  assign n508_o = n443_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n509_o = n446_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n510_o = n449_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n511_o = n452_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n512_o = n456_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n514_o = n461_o[2:0];
  /* upi41_core.vhd:394:3  */
  assign n515_o = n467_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n516_o = n473_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n517_o = n477_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n518_o = n480_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n519_o = n485_o[3:1];
  /* upi41_core.vhd:394:3  */
  assign n520_o = in_a_s[3:1];
  /* alu.vhd:200:5  */
  always @*
    case (n490_o)
      13'b1000000000000: n522_o = n520_o;
      13'b0100000000000: n522_o = n519_o;
      13'b0010000000000: n522_o = n518_o;
      13'b0001000000000: n522_o = n517_o;
      13'b0000100000000: n522_o = n516_o;
      13'b0000010000000: n522_o = n515_o;
      13'b0000001000000: n522_o = n514_o;
      13'b0000000100000: n522_o = 3'b000;
      13'b0000000010000: n522_o = n512_o;
      13'b0000000001000: n522_o = n511_o;
      13'b0000000000100: n522_o = n510_o;
      13'b0000000000010: n522_o = n509_o;
      13'b0000000000001: n522_o = n508_o;
      default: n522_o = 3'b000;
    endcase
  /* upi41_core.vhd:394:3  */
  assign n523_o = n443_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n524_o = n446_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n525_o = n449_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n526_o = n452_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n527_o = n456_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n529_o = n461_o[5:3];
  /* upi41_core.vhd:394:3  */
  assign n530_o = n467_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n531_o = n474_o[2:0];
  /* upi41_core.vhd:394:3  */
  assign n532_o = n477_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n533_o = n480_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n534_o = n485_o[6:4];
  /* upi41_core.vhd:394:3  */
  assign n535_o = in_a_s[6:4];
  /* alu.vhd:200:5  */
  always @*
    case (n490_o)
      13'b1000000000000: n537_o = n535_o;
      13'b0100000000000: n537_o = n534_o;
      13'b0010000000000: n537_o = n533_o;
      13'b0001000000000: n537_o = n532_o;
      13'b0000100000000: n537_o = n531_o;
      13'b0000010000000: n537_o = n530_o;
      13'b0000001000000: n537_o = n529_o;
      13'b0000000100000: n537_o = 3'b000;
      13'b0000000010000: n537_o = n527_o;
      13'b0000000001000: n537_o = n526_o;
      13'b0000000000100: n537_o = n525_o;
      13'b0000000000010: n537_o = n524_o;
      13'b0000000000001: n537_o = n523_o;
      default: n537_o = 3'b000;
    endcase
  /* upi41_core.vhd:394:3  */
  assign n538_o = n443_o[7];
  /* upi41_core.vhd:394:3  */
  assign n539_o = n446_o[7];
  /* upi41_core.vhd:394:3  */
  assign n540_o = n449_o[7];
  /* upi41_core.vhd:394:3  */
  assign n541_o = n452_o[7];
  /* upi41_core.vhd:394:3  */
  assign n542_o = n456_o[7];
  /* upi41_core.vhd:394:3  */
  assign n544_o = n461_o[6];
  /* upi41_core.vhd:394:3  */
  assign n545_o = n474_o[3];
  /* upi41_core.vhd:394:3  */
  assign n546_o = n477_o[7];
  /* upi41_core.vhd:394:3  */
  assign n547_o = n480_o[7];
  /* upi41_core.vhd:394:3  */
  assign n548_o = n485_o[7];
  /* upi41_core.vhd:394:3  */
  assign n549_o = in_a_s[7];
  /* alu.vhd:200:5  */
  always @*
    case (n490_o)
      13'b1000000000000: n551_o = n549_o;
      13'b0100000000000: n551_o = n548_o;
      13'b0010000000000: n551_o = n547_o;
      13'b0001000000000: n551_o = n546_o;
      13'b0000100000000: n551_o = n545_o;
      13'b0000010000000: n551_o = n470_o;
      13'b0000001000000: n551_o = n544_o;
      13'b0000000100000: n551_o = 1'b0;
      13'b0000000010000: n551_o = n542_o;
      13'b0000000001000: n551_o = n541_o;
      13'b0000000000100: n551_o = n540_o;
      13'b0000000000010: n551_o = n539_o;
      13'b0000000000001: n551_o = n538_o;
      default: n551_o = 1'b0;
    endcase
  /* alu.vhd:307:20  */
  assign n563_o = use_carry_i & carry_i;
  /* alu.vhd:307:5  */
  assign n566_o = n563_o ? 1'b1 : 1'b0;
  /* upi41_core.vhd:380:25  */
  assign n568_o = n567_o[8:1];
  /* alu.vhd:313:20  */
  assign n570_o = {1'b0, in_a_s};
  /* alu.vhd:314:20  */
  assign n572_o = {1'b0, in_b_s};
  /* upi41_core.vhd:356:5  */
  assign n575_o = n574_o[8:1];
  /* alu.vhd:317:7  */
  assign n577_o = alu_op_i == 4'b1001;
  /* alu.vhd:320:7  */
  assign n579_o = alu_op_i == 4'b1000;
  /* upi41_core.vhd:356:5  */
  assign n580_o = {n579_o, n577_o};
  /* upi41_core.vhd:356:5  */
  assign n582_o = n572_o[0];
  /* alu.vhd:316:5  */
  always @*
    case (n580_o)
      2'b10: n583_o = 1'b1;
      2'b01: n583_o = 1'b1;
      default: n583_o = n582_o;
    endcase
  /* upi41_core.vhd:356:5  */
  assign n585_o = n572_o[8:1];
  /* alu.vhd:316:5  */
  always @*
    case (n580_o)
      2'b10: n586_o = 8'b11111111;
      2'b01: n586_o = n575_o;
      default: n586_o = n585_o;
    endcase
  /* upi41_core.vhd:335:3  */
  assign n588_o = {n586_o, n583_o};
  /* alu.vhd:327:35  */
  assign n589_o = n570_o + n588_o;
  /* upi41_core.vhd:328:25  */
  assign n590_o = {n568_o, n566_o};
  /* alu.vhd:328:35  */
  assign n591_o = n589_o + n590_o;
  /* alu.vhd:334:32  */
  assign n592_o = in_a_s[4];
  /* alu.vhd:334:44  */
  assign n593_o = in_b_s[4];
  /* alu.vhd:334:36  */
  assign n594_o = {n592_o, n593_o};
  /* alu.vhd:339:20  */
  assign n595_o = n591_o[4];
  /* alu.vhd:339:9  */
  assign n598_o = n595_o ? 1'b1 : 1'b0;
  /* alu.vhd:338:7  */
  assign n600_o = n594_o == 2'b00;
  /* alu.vhd:338:17  */
  assign n602_o = n594_o == 2'b11;
  /* alu.vhd:338:17  */
  assign n603_o = n600_o | n602_o;
  /* alu.vhd:344:20  */
  assign n604_o = n591_o[4];
  /* alu.vhd:344:24  */
  assign n605_o = ~n604_o;
  /* alu.vhd:344:9  */
  assign n608_o = n605_o ? 1'b1 : 1'b0;
  /* alu.vhd:343:7  */
  assign n610_o = n594_o == 2'b01;
  /* alu.vhd:343:17  */
  assign n612_o = n594_o == 2'b10;
  /* alu.vhd:343:17  */
  assign n613_o = n610_o | n612_o;
  /* upi41_core.vhd:94:5  */
  assign n614_o = {n613_o, n603_o};
  /* alu.vhd:337:5  */
  always @*
    case (n614_o)
      2'b10: n616_o = n608_o;
      2'b01: n616_o = n598_o;
      default: n616_o = 1'b0;
    endcase
  /* alu.vhd:389:35  */
  assign n623_o = accu_shadow_q[7:4];
  /* alu.vhd:391:35  */
  assign n624_o = accu_shadow_q[3:0];
  /* alu.vhd:388:5  */
  assign n625_o = da_high_i ? n623_o : n624_o;
  /* alu.vhd:373:9  */
  assign n633_o = n625_o == 4'b1010;
  /* alu.vhd:373:21  */
  assign n635_o = n625_o == 4'b1011;
  /* alu.vhd:373:21  */
  assign n636_o = n633_o | n635_o;
  /* alu.vhd:374:21  */
  assign n638_o = n625_o == 4'b1100;
  /* alu.vhd:374:21  */
  assign n639_o = n636_o | n638_o;
  /* alu.vhd:375:21  */
  assign n641_o = n625_o == 4'b1101;
  /* alu.vhd:375:21  */
  assign n642_o = n639_o | n641_o;
  /* alu.vhd:376:21  */
  assign n644_o = n625_o == 4'b1110;
  /* alu.vhd:376:21  */
  assign n645_o = n642_o | n644_o;
  /* alu.vhd:377:21  */
  assign n647_o = n625_o == 4'b1111;
  /* alu.vhd:377:21  */
  assign n648_o = n645_o | n647_o;
  /* alu.vhd:372:7  */
  always @*
    case (n648_o)
      1'b1: n651_o = 1'b1;
      default: n651_o = 1'b0;
    endcase
  /* alu.vhd:412:13  */
  assign n654_o = read_alu_i ? data_s : 8'b11111111;
  /* alu.vhd:127:5  */
  assign n656_o = n429_o ? n421_o : accumulator_q;
  /* alu.vhd:127:5  */
  always @(posedge clk_i or posedge n413_o)
    if (n413_o)
      n657_q <= 8'b00000000;
    else
      n657_q <= n656_o;
  /* alu.vhd:127:5  */
  assign n658_o = en_clk_i ? n423_o : accu_shadow_q;
  /* alu.vhd:127:5  */
  always @(posedge clk_i or posedge n413_o)
    if (n413_o)
      n659_q <= 8'b00000000;
    else
      n659_q <= n658_o;
  /* alu.vhd:127:5  */
  assign n660_o = en_clk_i ? n428_o : temp_req_q;
  /* alu.vhd:127:5  */
  always @(posedge clk_i or posedge n413_o)
    if (n413_o)
      n661_q <= 8'b00000000;
    else
      n661_q <= n660_o;
  /* alu.vhd:122:5  */
  assign n662_o = {n551_o, n537_o, n522_o, n507_o};
endmodule

module upi41_core
  (input  xtal_i,
   input  xtal_en_i,
   input  reset_i,
   input  t0_i,
   input  cs_n_i,
   input  rd_n_i,
   input  a0_i,
   input  wr_n_i,
   input  [7:0] db_i,
   input  t1_i,
   input  [7:0] p2_i,
   input  [7:0] p1_i,
   input  clk_i,
   input  en_clk_i,
   input  [7:0] dmem_data_i,
   input  [7:0] pmem_data_i,
   output sync_o,
   output [7:0] db_o,
   output db_dir_o,
   output [7:0] p2_o,
   output p2l_low_imp_o,
   output p2h_low_imp_o,
   output [7:0] p1_o,
   output p1_low_imp_o,
   output prog_n_o,
   output xtal3_o,
   output [7:0] dmem_addr_o,
   output dmem_we_o,
   output [7:0] dmem_data_o,
   output [10:0] pmem_addr_o);
  wire [7:0] t48_data_s;
  wire xtal_en_s;
  wire en_clk_s;
  wire t0_s;
  wire t1_s;
  wire [7:0] alu_data_s;
  wire alu_write_accu_s;
  wire alu_write_shadow_s;
  wire alu_write_temp_reg_s;
  wire alu_read_alu_s;
  wire alu_carry_s;
  wire alu_aux_carry_s;
  wire [3:0] alu_op_s;
  wire alu_use_carry_s;
  wire alu_da_high_s;
  wire alu_da_overflow_s;
  wire alu_accu_low_s;
  wire alu_p06_temp_reg_s;
  wire alu_p60_temp_reg_s;
  wire bus_write_bus_s;
  wire bus_read_bus_s;
  wire [7:0] bus_data_s;
  wire bus_ibf_s;
  wire bus_obf_s;
  wire bus_int_n_s;
  wire bus_set_f1_s;
  wire bus_clear_f1_s;
  wire bus_ibf_int_s;
  wire bus_en_dma_s;
  wire bus_en_flags_s;
  wire bus_write_sts_s;
  wire bus_mint_ibf_n_s;
  wire bus_mint_obf_s;
  wire bus_dma_s;
  wire bus_drq_s;
  wire clk_multi_cycle_s;
  wire clk_assert_psen_s;
  wire clk_assert_prog_s;
  wire clk_assert_rd_s;
  wire clk_assert_wr_s;
  wire [2:0] clk_mstate_s;
  wire clk_second_cycle_s;
  wire prog_s;
  wire ale_s;
  wire xtal3_s;
  wire cnd_compute_take_s;
  wire [3:0] cnd_branch_cond_s;
  wire cnd_take_branch_s;
  wire [2:0] cnd_comp_value_s;
  wire cnd_f1_s;
  wire cnd_tf_s;
  wire dm_write_dmem_addr_s;
  wire dm_write_dmem_s;
  wire dm_read_dmem_s;
  wire [1:0] dm_addr_type_s;
  wire [7:0] dm_data_s;
  wire [7:0] dec_data_s;
  wire p1_write_p1_s;
  wire p1_read_p1_s;
  wire p1_read_reg_s;
  wire [7:0] p1_data_s;
  wire [7:0] p2_s;
  wire p26_s;
  wire p2_write_p2_s;
  wire p2_write_exp_s;
  wire p2_read_p2_s;
  wire p2_read_reg_s;
  wire p2_read_exp_s;
  wire p2_output_pch_s;
  wire [7:0] p2_data_s;
  wire pm_write_pcl_s;
  wire pm_read_pcl_s;
  wire pm_write_pch_s;
  wire pm_read_pch_s;
  wire pm_read_pmem_s;
  wire pm_inc_pc_s;
  wire pm_write_pmem_addr_s;
  wire [7:0] pm_data_s;
  wire [1:0] pm_addr_type_s;
  wire [11:0] pmem_addr_s;
  wire psw_read_psw_s;
  wire psw_read_sp_s;
  wire psw_write_psw_s;
  wire psw_write_sp_s;
  wire psw_carry_s;
  wire psw_aux_carry_s;
  wire psw_f0_s;
  wire psw_bs_s;
  wire psw_special_data_s;
  wire psw_inc_stackp_s;
  wire psw_dec_stackp_s;
  wire psw_write_carry_s;
  wire psw_write_aux_carry_s;
  wire psw_write_f0_s;
  wire psw_write_bs_s;
  wire [7:0] psw_data_s;
  wire tim_overflow_s;
  wire tim_of_s;
  wire tim_read_timer_s;
  wire tim_write_timer_s;
  wire tim_start_t_s;
  wire tim_start_cnt_s;
  wire tim_stop_tcnt_s;
  wire [7:0] tim_data_s;
  wire gnd_s;
  localparam n14_o = 1'b0;
  wire n23_o;
  wire n31_o;
  wire [7:0] alu_b_n32;
  wire alu_b_n33;
  wire alu_b_n34;
  wire alu_b_n35;
  wire [7:0] alu_b_data_o;
  wire alu_b_carry_o;
  wire alu_b_aux_carry_o;
  wire alu_b_da_overflow_o;
  wire [7:0] bus_mux_b_n44;
  wire [7:0] bus_mux_b_data_o;
  wire clock_ctrl_b_n47;
  wire [2:0] clock_ctrl_b_n49;
  wire clock_ctrl_b_n50;
  wire clock_ctrl_b_n51;
  wire clock_ctrl_b_n53;
  wire clock_ctrl_b_xtal3_o;
  wire clock_ctrl_b_t0_o;
  wire [2:0] clock_ctrl_b_mstate_o;
  wire clock_ctrl_b_second_cycle_o;
  wire clock_ctrl_b_ale_o;
  wire clock_ctrl_b_psen_o;
  wire clock_ctrl_b_prog_o;
  wire clock_ctrl_b_rd_o;
  wire clock_ctrl_b_wr_o;
  wire cond_branch_b_n70;
  wire cond_branch_b_take_branch_o;
  wire [7:0] db_bus_b_n73;
  wire db_bus_b_n74;
  wire db_bus_b_n75;
  wire db_bus_b_n76;
  wire db_bus_b_n77;
  wire db_bus_b_n78;
  wire db_bus_b_n79;
  wire db_bus_b_n80;
  wire db_bus_b_n81;
  wire db_bus_b_n82;
  wire n83_o;
  wire [7:0] db_bus_b_n84;
  wire db_bus_b_n85;
  wire [7:0] db_bus_b_data_o;
  wire db_bus_b_set_f1_o;
  wire db_bus_b_clear_f1_o;
  wire db_bus_b_ibf_o;
  wire db_bus_b_obf_o;
  wire db_bus_b_int_n_o;
  wire db_bus_b_mint_ibf_n_o;
  wire db_bus_b_mint_obf_o;
  wire db_bus_b_dma_o;
  wire db_bus_b_drq_o;
  wire [7:0] db_bus_b_db_o;
  wire db_bus_b_db_dir_o;
  wire [7:0] decoder_b_n111;
  wire decoder_b_n112;
  wire decoder_b_n113;
  wire decoder_b_n114;
  wire decoder_b_n115;
  wire decoder_b_n116;
  wire decoder_b_n117;
  wire decoder_b_n118;
  wire decoder_b_n119;
  wire decoder_b_n120;
  wire decoder_b_n121;
  wire decoder_b_n122;
  wire decoder_b_n123;
  wire decoder_b_n124;
  wire decoder_b_n125;
  wire decoder_b_n126;
  wire decoder_b_n127;
  wire decoder_b_n128;
  wire decoder_b_n129;
  wire decoder_b_n130;
  wire decoder_b_n131;
  wire decoder_b_n132;
  wire decoder_b_n133;
  wire decoder_b_n134;
  wire decoder_b_n135;
  wire decoder_b_n136;
  wire decoder_b_n137;
  wire decoder_b_n138;
  wire [3:0] decoder_b_n139;
  wire decoder_b_n140;
  wire decoder_b_n141;
  wire decoder_b_n142;
  wire decoder_b_n143;
  wire decoder_b_n144;
  wire decoder_b_n147;
  wire decoder_b_n148;
  wire decoder_b_n149;
  wire decoder_b_n150;
  wire decoder_b_n151;
  wire decoder_b_n152;
  wire [3:0] decoder_b_n153;
  wire [2:0] decoder_b_n154;
  wire decoder_b_n155;
  wire decoder_b_n156;
  wire [1:0] decoder_b_n157;
  wire decoder_b_n158;
  wire decoder_b_n159;
  wire decoder_b_n160;
  wire decoder_b_n161;
  wire decoder_b_n162;
  wire decoder_b_n163;
  wire decoder_b_n164;
  wire decoder_b_n165;
  wire decoder_b_n166;
  wire decoder_b_n167;
  wire decoder_b_n168;
  wire [1:0] decoder_b_n169;
  wire decoder_b_n170;
  wire decoder_b_n171;
  wire decoder_b_n172;
  wire decoder_b_n173;
  wire decoder_b_n174;
  wire decoder_b_n175;
  wire decoder_b_n176;
  wire decoder_b_t0_dir_o;
  wire [7:0] decoder_b_data_o;
  wire decoder_b_alu_write_accu_o;
  wire decoder_b_alu_write_shadow_o;
  wire decoder_b_alu_write_temp_reg_o;
  wire decoder_b_alu_read_alu_o;
  wire decoder_b_bus_write_bus_o;
  wire decoder_b_bus_read_bus_o;
  wire decoder_b_bus_ibf_int_o;
  wire decoder_b_bus_en_dma_o;
  wire decoder_b_bus_en_flags_o;
  wire decoder_b_bus_write_sts_o;
  wire decoder_b_dm_write_dmem_addr_o;
  wire decoder_b_dm_write_dmem_o;
  wire decoder_b_dm_read_dmem_o;
  wire decoder_b_p1_write_p1_o;
  wire decoder_b_p1_read_p1_o;
  wire decoder_b_p2_write_p2_o;
  wire decoder_b_p2_write_exp_o;
  wire decoder_b_p2_read_p2_o;
  wire decoder_b_p2_read_exp_o;
  wire decoder_b_pm_write_pcl_o;
  wire decoder_b_pm_read_pcl_o;
  wire decoder_b_pm_write_pch_o;
  wire decoder_b_pm_read_pch_o;
  wire decoder_b_pm_read_pmem_o;
  wire decoder_b_psw_read_psw_o;
  wire decoder_b_psw_read_sp_o;
  wire decoder_b_psw_write_psw_o;
  wire decoder_b_psw_write_sp_o;
  wire [3:0] decoder_b_alu_op_o;
  wire decoder_b_alu_use_carry_o;
  wire decoder_b_alu_da_high_o;
  wire decoder_b_alu_accu_low_o;
  wire decoder_b_alu_p06_temp_reg_o;
  wire decoder_b_alu_p60_temp_reg_o;
  wire decoder_b_bus_output_pcl_o;
  wire decoder_b_bus_bidir_bus_o;
  wire decoder_b_clk_multi_cycle_o;
  wire decoder_b_clk_assert_psen_o;
  wire decoder_b_clk_assert_prog_o;
  wire decoder_b_clk_assert_rd_o;
  wire decoder_b_clk_assert_wr_o;
  wire decoder_b_cnd_compute_take_o;
  wire [3:0] decoder_b_cnd_branch_cond_o;
  wire [2:0] decoder_b_cnd_comp_value_o;
  wire decoder_b_cnd_f1_o;
  wire decoder_b_cnd_tf_o;
  wire [1:0] decoder_b_dm_addr_type_o;
  wire decoder_b_p1_read_reg_o;
  wire decoder_b_p2_read_reg_o;
  wire decoder_b_p2_output_pch_o;
  wire decoder_b_pm_inc_pc_o;
  wire decoder_b_pm_write_pmem_addr_o;
  wire [1:0] decoder_b_pm_addr_type_o;
  wire decoder_b_psw_special_data_o;
  wire decoder_b_psw_inc_stackp_o;
  wire decoder_b_psw_dec_stackp_o;
  wire decoder_b_psw_write_carry_o;
  wire decoder_b_psw_write_aux_carry_o;
  wire decoder_b_psw_write_f0_o;
  wire decoder_b_psw_write_bs_o;
  wire decoder_b_tim_read_timer_o;
  wire decoder_b_tim_write_timer_o;
  wire decoder_b_tim_start_t_o;
  wire decoder_b_tim_start_cnt_o;
  wire decoder_b_tim_stop_tcnt_o;
  wire [7:0] dmem_ctrl_b_n308;
  wire [7:0] dmem_ctrl_b_n309;
  wire dmem_ctrl_b_n310;
  wire [7:0] dmem_ctrl_b_n311;
  wire [7:0] dmem_ctrl_b_data_o;
  wire [7:0] dmem_ctrl_b_dmem_addr_o;
  wire dmem_ctrl_b_dmem_we_o;
  wire [7:0] dmem_ctrl_b_dmem_data_o;
  wire [7:0] timer_b_n320;
  wire timer_b_n321;
  wire [7:0] timer_b_data_o;
  wire timer_b_overflow_o;
  wire n333_o;
  wire [7:0] p1_b_n334;
  wire [7:0] p1_b_n335;
  wire p1_b_n336;
  wire [7:0] p1_b_data_o;
  wire [7:0] p1_b_p1_o;
  wire p1_b_p1_low_imp_o;
  wire [7:0] p2_b_n343;
  wire [3:0] n344_o;
  wire [7:0] p2_b_n345;
  wire p2_b_n346;
  wire p2_b_n347;
  wire [7:0] p2_b_data_o;
  wire [7:0] p2_b_p2_o;
  wire p2_b_p2l_low_imp_o;
  wire p2_b_p2h_low_imp_o;
  wire n356_o;
  wire n357_o;
  wire n358_o;
  wire n359_o;
  wire [1:0] n360_o;
  wire n361_o;
  wire n362_o;
  wire [2:0] n363_o;
  wire n364_o;
  wire n365_o;
  wire [3:0] n366_o;
  wire [3:0] n367_o;
  wire [7:0] n368_o;
  wire [7:0] pmem_ctrl_b_n369;
  wire [11:0] pmem_ctrl_b_n370;
  wire [7:0] pmem_ctrl_b_data_o;
  wire [11:0] pmem_ctrl_b_pmem_addr_o;
  wire [7:0] psw_b_n375;
  wire psw_b_n376;
  wire psw_b_n377;
  wire psw_b_n378;
  wire psw_b_n379;
  wire [7:0] psw_b_data_o;
  wire psw_b_carry_o;
  wire psw_b_aux_carry_o;
  wire psw_b_f0_o;
  wire psw_b_bs_o;
  wire n391_o;
  wire n398_o;
  wire n406_o;
  wire [10:0] n407_o;
  assign sync_o = n14_o;
  assign db_o = db_bus_b_n84;
  assign db_dir_o = db_bus_b_n85;
  assign p2_o = n368_o;
  assign p2l_low_imp_o = p2_b_n346;
  assign p2h_low_imp_o = p2_b_n347;
  assign p1_o = p1_b_n335;
  assign p1_low_imp_o = p1_b_n336;
  assign prog_n_o = n398_o;
  assign xtal3_o = n406_o;
  assign dmem_addr_o = dmem_ctrl_b_n309;
  assign dmem_we_o = dmem_ctrl_b_n310;
  assign dmem_data_o = dmem_ctrl_b_n311;
  assign pmem_addr_o = n407_o;
  /* upi41_core.vhd:125:10  */
  assign t48_data_s = bus_mux_b_n44; // (signal)
  /* upi41_core.vhd:127:10  */
  assign xtal_en_s = n23_o; // (signal)
  /* upi41_core.vhd:128:10  */
  assign en_clk_s = n31_o; // (signal)
  /* upi41_core.vhd:130:10  */
  assign t0_s = t0_i; // (signal)
  /* upi41_core.vhd:130:16  */
  assign t1_s = t1_i; // (signal)
  /* upi41_core.vhd:133:10  */
  assign alu_data_s = alu_b_n32; // (signal)
  /* upi41_core.vhd:134:10  */
  assign alu_write_accu_s = decoder_b_n112; // (signal)
  /* upi41_core.vhd:135:10  */
  assign alu_write_shadow_s = decoder_b_n113; // (signal)
  /* upi41_core.vhd:136:10  */
  assign alu_write_temp_reg_s = decoder_b_n114; // (signal)
  /* upi41_core.vhd:137:10  */
  assign alu_read_alu_s = decoder_b_n115; // (signal)
  /* upi41_core.vhd:138:10  */
  assign alu_carry_s = alu_b_n33; // (signal)
  /* upi41_core.vhd:139:10  */
  assign alu_aux_carry_s = alu_b_n34; // (signal)
  /* upi41_core.vhd:140:10  */
  assign alu_op_s = decoder_b_n139; // (signal)
  /* upi41_core.vhd:141:10  */
  assign alu_use_carry_s = decoder_b_n144; // (signal)
  /* upi41_core.vhd:142:10  */
  assign alu_da_high_s = decoder_b_n140; // (signal)
  /* upi41_core.vhd:143:10  */
  assign alu_da_overflow_s = alu_b_n35; // (signal)
  /* upi41_core.vhd:144:10  */
  assign alu_accu_low_s = decoder_b_n141; // (signal)
  /* upi41_core.vhd:145:10  */
  assign alu_p06_temp_reg_s = decoder_b_n142; // (signal)
  /* upi41_core.vhd:146:10  */
  assign alu_p60_temp_reg_s = decoder_b_n143; // (signal)
  /* upi41_core.vhd:149:10  */
  assign bus_write_bus_s = decoder_b_n116; // (signal)
  /* upi41_core.vhd:150:10  */
  assign bus_read_bus_s = decoder_b_n117; // (signal)
  /* upi41_core.vhd:151:10  */
  assign bus_data_s = db_bus_b_n73; // (signal)
  /* upi41_core.vhd:153:10  */
  assign bus_ibf_s = db_bus_b_n76; // (signal)
  /* upi41_core.vhd:154:10  */
  assign bus_obf_s = db_bus_b_n77; // (signal)
  /* upi41_core.vhd:155:10  */
  assign bus_int_n_s = db_bus_b_n78; // (signal)
  /* upi41_core.vhd:156:10  */
  assign bus_set_f1_s = db_bus_b_n74; // (signal)
  /* upi41_core.vhd:157:10  */
  assign bus_clear_f1_s = db_bus_b_n75; // (signal)
  /* upi41_core.vhd:158:10  */
  assign bus_ibf_int_s = decoder_b_n118; // (signal)
  /* upi41_core.vhd:159:10  */
  assign bus_en_dma_s = decoder_b_n119; // (signal)
  /* upi41_core.vhd:160:10  */
  assign bus_en_flags_s = decoder_b_n120; // (signal)
  /* upi41_core.vhd:161:10  */
  assign bus_write_sts_s = decoder_b_n121; // (signal)
  /* upi41_core.vhd:162:10  */
  assign bus_mint_ibf_n_s = db_bus_b_n79; // (signal)
  /* upi41_core.vhd:163:10  */
  assign bus_mint_obf_s = db_bus_b_n80; // (signal)
  /* upi41_core.vhd:164:10  */
  assign bus_dma_s = db_bus_b_n81; // (signal)
  /* upi41_core.vhd:165:10  */
  assign bus_drq_s = db_bus_b_n82; // (signal)
  /* upi41_core.vhd:168:10  */
  assign clk_multi_cycle_s = decoder_b_n147; // (signal)
  /* upi41_core.vhd:169:10  */
  assign clk_assert_psen_s = decoder_b_n148; // (signal)
  /* upi41_core.vhd:170:10  */
  assign clk_assert_prog_s = decoder_b_n149; // (signal)
  /* upi41_core.vhd:171:10  */
  assign clk_assert_rd_s = decoder_b_n150; // (signal)
  /* upi41_core.vhd:172:10  */
  assign clk_assert_wr_s = decoder_b_n151; // (signal)
  /* upi41_core.vhd:173:10  */
  assign clk_mstate_s = clock_ctrl_b_n49; // (signal)
  /* upi41_core.vhd:174:10  */
  assign clk_second_cycle_s = clock_ctrl_b_n50; // (signal)
  /* upi41_core.vhd:175:10  */
  assign prog_s = clock_ctrl_b_n53; // (signal)
  /* upi41_core.vhd:176:10  */
  assign ale_s = clock_ctrl_b_n51; // (signal)
  /* upi41_core.vhd:177:10  */
  assign xtal3_s = clock_ctrl_b_n47; // (signal)
  /* upi41_core.vhd:180:10  */
  assign cnd_compute_take_s = decoder_b_n152; // (signal)
  /* upi41_core.vhd:181:10  */
  assign cnd_branch_cond_s = decoder_b_n153; // (signal)
  /* upi41_core.vhd:182:10  */
  assign cnd_take_branch_s = cond_branch_b_n70; // (signal)
  /* upi41_core.vhd:183:10  */
  assign cnd_comp_value_s = decoder_b_n154; // (signal)
  /* upi41_core.vhd:184:10  */
  assign cnd_f1_s = decoder_b_n155; // (signal)
  /* upi41_core.vhd:185:10  */
  assign cnd_tf_s = decoder_b_n156; // (signal)
  /* upi41_core.vhd:188:10  */
  assign dm_write_dmem_addr_s = decoder_b_n122; // (signal)
  /* upi41_core.vhd:189:10  */
  assign dm_write_dmem_s = decoder_b_n123; // (signal)
  /* upi41_core.vhd:190:10  */
  assign dm_read_dmem_s = decoder_b_n124; // (signal)
  /* upi41_core.vhd:191:10  */
  assign dm_addr_type_s = decoder_b_n157; // (signal)
  /* upi41_core.vhd:192:10  */
  assign dm_data_s = dmem_ctrl_b_n308; // (signal)
  /* upi41_core.vhd:195:10  */
  assign dec_data_s = decoder_b_n111; // (signal)
  /* upi41_core.vhd:198:10  */
  assign p1_write_p1_s = decoder_b_n125; // (signal)
  /* upi41_core.vhd:199:10  */
  assign p1_read_p1_s = decoder_b_n126; // (signal)
  /* upi41_core.vhd:200:10  */
  assign p1_read_reg_s = decoder_b_n163; // (signal)
  /* upi41_core.vhd:201:10  */
  assign p1_data_s = p1_b_n334; // (signal)
  /* upi41_core.vhd:204:10  */
  assign p2_s = p2_b_n345; // (signal)
  /* upi41_core.vhd:205:10  */
  assign p26_s = n358_o; // (signal)
  /* upi41_core.vhd:206:10  */
  assign p2_write_p2_s = decoder_b_n127; // (signal)
  /* upi41_core.vhd:207:10  */
  assign p2_write_exp_s = decoder_b_n128; // (signal)
  /* upi41_core.vhd:208:10  */
  assign p2_read_p2_s = decoder_b_n129; // (signal)
  /* upi41_core.vhd:209:10  */
  assign p2_read_reg_s = decoder_b_n164; // (signal)
  /* upi41_core.vhd:210:10  */
  assign p2_read_exp_s = decoder_b_n165; // (signal)
  /* upi41_core.vhd:211:10  */
  assign p2_output_pch_s = decoder_b_n166; // (signal)
  /* upi41_core.vhd:212:10  */
  assign p2_data_s = p2_b_n343; // (signal)
  /* upi41_core.vhd:215:10  */
  assign pm_write_pcl_s = decoder_b_n130; // (signal)
  /* upi41_core.vhd:216:10  */
  assign pm_read_pcl_s = decoder_b_n131; // (signal)
  /* upi41_core.vhd:217:10  */
  assign pm_write_pch_s = decoder_b_n132; // (signal)
  /* upi41_core.vhd:218:10  */
  assign pm_read_pch_s = decoder_b_n133; // (signal)
  /* upi41_core.vhd:219:10  */
  assign pm_read_pmem_s = decoder_b_n134; // (signal)
  /* upi41_core.vhd:220:10  */
  assign pm_inc_pc_s = decoder_b_n167; // (signal)
  /* upi41_core.vhd:221:10  */
  assign pm_write_pmem_addr_s = decoder_b_n168; // (signal)
  /* upi41_core.vhd:222:10  */
  assign pm_data_s = pmem_ctrl_b_n369; // (signal)
  /* upi41_core.vhd:223:10  */
  assign pm_addr_type_s = decoder_b_n169; // (signal)
  /* upi41_core.vhd:224:10  */
  assign pmem_addr_s = pmem_ctrl_b_n370; // (signal)
  /* upi41_core.vhd:227:10  */
  assign psw_read_psw_s = decoder_b_n135; // (signal)
  /* upi41_core.vhd:228:10  */
  assign psw_read_sp_s = decoder_b_n136; // (signal)
  /* upi41_core.vhd:229:10  */
  assign psw_write_psw_s = decoder_b_n137; // (signal)
  /* upi41_core.vhd:230:10  */
  assign psw_write_sp_s = decoder_b_n138; // (signal)
  /* upi41_core.vhd:231:10  */
  assign psw_carry_s = psw_b_n376; // (signal)
  /* upi41_core.vhd:232:10  */
  assign psw_aux_carry_s = psw_b_n377; // (signal)
  /* upi41_core.vhd:233:10  */
  assign psw_f0_s = psw_b_n378; // (signal)
  /* upi41_core.vhd:234:10  */
  assign psw_bs_s = psw_b_n379; // (signal)
  /* upi41_core.vhd:235:10  */
  assign psw_special_data_s = decoder_b_n170; // (signal)
  /* upi41_core.vhd:236:10  */
  assign psw_inc_stackp_s = decoder_b_n171; // (signal)
  /* upi41_core.vhd:237:10  */
  assign psw_dec_stackp_s = decoder_b_n172; // (signal)
  /* upi41_core.vhd:238:10  */
  assign psw_write_carry_s = decoder_b_n173; // (signal)
  /* upi41_core.vhd:239:10  */
  assign psw_write_aux_carry_s = decoder_b_n174; // (signal)
  /* upi41_core.vhd:240:10  */
  assign psw_write_f0_s = decoder_b_n175; // (signal)
  /* upi41_core.vhd:241:10  */
  assign psw_write_bs_s = decoder_b_n176; // (signal)
  /* upi41_core.vhd:242:10  */
  assign psw_data_s = psw_b_n375; // (signal)
  /* upi41_core.vhd:245:10  */
  assign tim_overflow_s = n333_o; // (signal)
  /* upi41_core.vhd:246:10  */
  assign tim_of_s = timer_b_n321; // (signal)
  /* upi41_core.vhd:247:10  */
  assign tim_read_timer_s = decoder_b_n158; // (signal)
  /* upi41_core.vhd:248:10  */
  assign tim_write_timer_s = decoder_b_n159; // (signal)
  /* upi41_core.vhd:249:10  */
  assign tim_start_t_s = decoder_b_n160; // (signal)
  /* upi41_core.vhd:250:10  */
  assign tim_start_cnt_s = decoder_b_n161; // (signal)
  /* upi41_core.vhd:251:10  */
  assign tim_stop_tcnt_s = decoder_b_n162; // (signal)
  /* upi41_core.vhd:252:10  */
  assign tim_data_s = timer_b_n320; // (signal)
  /* upi41_core.vhd:254:10  */
  assign gnd_s = 1'b0; // (signal)
  /* t48_pack-p.vhd:75:5  */
  assign n23_o = xtal_en_i ? 1'b1 : 1'b0;
  /* t48_pack-p.vhd:75:5  */
  assign n31_o = en_clk_i ? 1'b1 : 1'b0;
  /* upi41_core.vhd:278:29  */
  assign alu_b_n32 = alu_b_data_o; // (signal)
  /* upi41_core.vhd:284:29  */
  assign alu_b_n33 = alu_b_carry_o; // (signal)
  /* upi41_core.vhd:285:29  */
  assign alu_b_n34 = alu_b_aux_carry_o; // (signal)
  /* upi41_core.vhd:289:29  */
  assign alu_b_n35 = alu_b_da_overflow_o; // (signal)
  /* upi41_core.vhd:272:3  */
  t48_alu alu_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_accu_i(alu_write_accu_s),
    .write_shadow_i(alu_write_shadow_s),
    .write_temp_reg_i(alu_write_temp_reg_s),
    .read_alu_i(alu_read_alu_s),
    .carry_i(psw_carry_s),
    .alu_op_i(alu_op_s),
    .use_carry_i(alu_use_carry_s),
    .da_high_i(alu_da_high_s),
    .accu_low_i(alu_accu_low_s),
    .p06_temp_reg_i(alu_p06_temp_reg_s),
    .p60_temp_reg_i(alu_p60_temp_reg_s),
    .data_o(alu_b_data_o),
    .carry_o(alu_b_carry_o),
    .aux_carry_o(alu_b_aux_carry_o),
    .da_overflow_o(alu_b_da_overflow_o));
  /* upi41_core.vhd:306:21  */
  assign bus_mux_b_n44 = bus_mux_b_data_o; // (signal)
  /* upi41_core.vhd:295:3  */
  t48_bus_mux bus_mux_b (
    .alu_data_i(alu_data_s),
    .bus_data_i(bus_data_s),
    .dec_data_i(dec_data_s),
    .dm_data_i(dm_data_s),
    .pm_data_i(pm_data_s),
    .p1_data_i(p1_data_s),
    .p2_data_i(p2_data_s),
    .psw_data_i(psw_data_s),
    .tim_data_i(tim_data_s),
    .data_o(bus_mux_b_data_o));
  /* upi41_core.vhd:319:25  */
  assign clock_ctrl_b_n47 = clock_ctrl_b_xtal3_o; // (signal)
  /* upi41_core.vhd:326:25  */
  assign clock_ctrl_b_n49 = clock_ctrl_b_mstate_o; // (signal)
  /* upi41_core.vhd:327:25  */
  assign clock_ctrl_b_n50 = clock_ctrl_b_second_cycle_o; // (signal)
  /* upi41_core.vhd:328:25  */
  assign clock_ctrl_b_n51 = clock_ctrl_b_ale_o; // (signal)
  /* upi41_core.vhd:330:25  */
  assign clock_ctrl_b_n53 = clock_ctrl_b_prog_o; // (signal)
  /* upi41_core.vhd:309:3  */
  t48_clock_ctrl_1 clock_ctrl_b (
    .clk_i(clk_i),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_s),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .multi_cycle_i(clk_multi_cycle_s),
    .assert_psen_i(clk_assert_psen_s),
    .assert_prog_i(clk_assert_prog_s),
    .assert_rd_i(clk_assert_rd_s),
    .assert_wr_i(clk_assert_wr_s),
    .xtal3_o(clock_ctrl_b_xtal3_o),
    .t0_o(),
    .mstate_o(clock_ctrl_b_mstate_o),
    .second_cycle_o(clock_ctrl_b_second_cycle_o),
    .ale_o(clock_ctrl_b_ale_o),
    .psen_o(),
    .prog_o(clock_ctrl_b_prog_o),
    .rd_o(),
    .wr_o());
  /* upi41_core.vhd:342:25  */
  assign cond_branch_b_n70 = cond_branch_b_take_branch_o; // (signal)
  /* upi41_core.vhd:335:3  */
  t48_cond_branch cond_branch_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .compute_take_i(cnd_compute_take_s),
    .branch_cond_i(cnd_branch_cond_s),
    .accu_i(alu_data_s),
    .t0_i(t0_s),
    .t1_i(t1_s),
    .int_n_i(bus_int_n_s),
    .f0_i(psw_f0_s),
    .f1_i(cnd_f1_s),
    .tf_i(cnd_tf_s),
    .carry_i(psw_carry_s),
    .ibf_i(bus_ibf_s),
    .obf_i(bus_obf_s),
    .comp_value_i(cnd_comp_value_s),
    .take_branch_o(cond_branch_b_take_branch_o));
  /* upi41_core.vhd:365:25  */
  assign db_bus_b_n73 = db_bus_b_data_o; // (signal)
  /* upi41_core.vhd:369:25  */
  assign db_bus_b_n74 = db_bus_b_set_f1_o; // (signal)
  /* upi41_core.vhd:370:25  */
  assign db_bus_b_n75 = db_bus_b_clear_f1_o; // (signal)
  /* upi41_core.vhd:373:25  */
  assign db_bus_b_n76 = db_bus_b_ibf_o; // (signal)
  /* upi41_core.vhd:374:25  */
  assign db_bus_b_n77 = db_bus_b_obf_o; // (signal)
  /* upi41_core.vhd:375:25  */
  assign db_bus_b_n78 = db_bus_b_int_n_o; // (signal)
  /* upi41_core.vhd:380:25  */
  assign db_bus_b_n79 = db_bus_b_mint_ibf_n_o; // (signal)
  /* upi41_core.vhd:381:25  */
  assign db_bus_b_n80 = db_bus_b_mint_obf_o; // (signal)
  /* upi41_core.vhd:382:25  */
  assign db_bus_b_n81 = db_bus_b_dma_o; // (signal)
  /* upi41_core.vhd:383:25  */
  assign db_bus_b_n82 = db_bus_b_drq_o; // (signal)
  /* upi41_core.vhd:384:29  */
  assign n83_o = p2_i[7];
  /* upi41_core.vhd:390:25  */
  assign db_bus_b_n84 = db_bus_b_db_o; // (signal)
  /* upi41_core.vhd:391:25  */
  assign db_bus_b_n85 = db_bus_b_db_dir_o; // (signal)
  /* upi41_core.vhd:356:5  */
  upi41_db_bus_1 db_bus_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_bus_i(bus_write_bus_s),
    .read_bus_i(bus_read_bus_s),
    .write_sts_i(bus_write_sts_s),
    .f0_i(psw_f0_s),
    .f1_i(cnd_f1_s),
    .ibf_int_i(bus_ibf_int_s),
    .en_dma_i(bus_en_dma_s),
    .en_flags_i(bus_en_flags_s),
    .write_p2_i(p2_write_p2_s),
    .dack_n_i(n83_o),
    .a0_i(a0_i),
    .cs_n_i(cs_n_i),
    .rd_n_i(rd_n_i),
    .wr_n_i(wr_n_i),
    .db_i(db_i),
    .data_o(db_bus_b_data_o),
    .set_f1_o(db_bus_b_set_f1_o),
    .clear_f1_o(db_bus_b_clear_f1_o),
    .ibf_o(db_bus_b_ibf_o),
    .obf_o(db_bus_b_obf_o),
    .int_n_o(db_bus_b_int_n_o),
    .mint_ibf_n_o(db_bus_b_mint_ibf_n_o),
    .mint_obf_o(db_bus_b_mint_obf_o),
    .dma_o(db_bus_b_dma_o),
    .drq_o(db_bus_b_drq_o),
    .db_o(db_bus_b_db_o),
    .db_dir_o(db_bus_b_db_dir_o));
  /* upi41_core.vhd:411:33  */
  assign decoder_b_n111 = decoder_b_data_o; // (signal)
  /* upi41_core.vhd:412:33  */
  assign decoder_b_n112 = decoder_b_alu_write_accu_o; // (signal)
  /* upi41_core.vhd:413:33  */
  assign decoder_b_n113 = decoder_b_alu_write_shadow_o; // (signal)
  /* upi41_core.vhd:414:33  */
  assign decoder_b_n114 = decoder_b_alu_write_temp_reg_o; // (signal)
  /* upi41_core.vhd:415:33  */
  assign decoder_b_n115 = decoder_b_alu_read_alu_o; // (signal)
  /* upi41_core.vhd:416:33  */
  assign decoder_b_n116 = decoder_b_bus_write_bus_o; // (signal)
  /* upi41_core.vhd:417:33  */
  assign decoder_b_n117 = decoder_b_bus_read_bus_o; // (signal)
  /* upi41_core.vhd:420:33  */
  assign decoder_b_n118 = decoder_b_bus_ibf_int_o; // (signal)
  /* upi41_core.vhd:421:33  */
  assign decoder_b_n119 = decoder_b_bus_en_dma_o; // (signal)
  /* upi41_core.vhd:422:33  */
  assign decoder_b_n120 = decoder_b_bus_en_flags_o; // (signal)
  /* upi41_core.vhd:423:33  */
  assign decoder_b_n121 = decoder_b_bus_write_sts_o; // (signal)
  /* upi41_core.vhd:424:33  */
  assign decoder_b_n122 = decoder_b_dm_write_dmem_addr_o; // (signal)
  /* upi41_core.vhd:425:33  */
  assign decoder_b_n123 = decoder_b_dm_write_dmem_o; // (signal)
  /* upi41_core.vhd:426:33  */
  assign decoder_b_n124 = decoder_b_dm_read_dmem_o; // (signal)
  /* upi41_core.vhd:427:33  */
  assign decoder_b_n125 = decoder_b_p1_write_p1_o; // (signal)
  /* upi41_core.vhd:428:33  */
  assign decoder_b_n126 = decoder_b_p1_read_p1_o; // (signal)
  /* upi41_core.vhd:430:33  */
  assign decoder_b_n127 = decoder_b_p2_write_p2_o; // (signal)
  /* upi41_core.vhd:431:33  */
  assign decoder_b_n128 = decoder_b_p2_write_exp_o; // (signal)
  /* upi41_core.vhd:432:33  */
  assign decoder_b_n129 = decoder_b_p2_read_p2_o; // (signal)
  /* upi41_core.vhd:429:33  */
  assign decoder_b_n130 = decoder_b_pm_write_pcl_o; // (signal)
  /* upi41_core.vhd:433:33  */
  assign decoder_b_n131 = decoder_b_pm_read_pcl_o; // (signal)
  /* upi41_core.vhd:434:33  */
  assign decoder_b_n132 = decoder_b_pm_write_pch_o; // (signal)
  /* upi41_core.vhd:435:33  */
  assign decoder_b_n133 = decoder_b_pm_read_pch_o; // (signal)
  /* upi41_core.vhd:436:33  */
  assign decoder_b_n134 = decoder_b_pm_read_pmem_o; // (signal)
  /* upi41_core.vhd:437:33  */
  assign decoder_b_n135 = decoder_b_psw_read_psw_o; // (signal)
  /* upi41_core.vhd:438:33  */
  assign decoder_b_n136 = decoder_b_psw_read_sp_o; // (signal)
  /* upi41_core.vhd:439:33  */
  assign decoder_b_n137 = decoder_b_psw_write_psw_o; // (signal)
  /* upi41_core.vhd:440:33  */
  assign decoder_b_n138 = decoder_b_psw_write_sp_o; // (signal)
  /* upi41_core.vhd:442:33  */
  assign decoder_b_n139 = decoder_b_alu_op_o; // (signal)
  /* upi41_core.vhd:444:33  */
  assign decoder_b_n140 = decoder_b_alu_da_high_o; // (signal)
  /* upi41_core.vhd:446:33  */
  assign decoder_b_n141 = decoder_b_alu_accu_low_o; // (signal)
  /* upi41_core.vhd:447:33  */
  assign decoder_b_n142 = decoder_b_alu_p06_temp_reg_o; // (signal)
  /* upi41_core.vhd:448:33  */
  assign decoder_b_n143 = decoder_b_alu_p60_temp_reg_o; // (signal)
  /* upi41_core.vhd:443:33  */
  assign decoder_b_n144 = decoder_b_alu_use_carry_o; // (signal)
  /* upi41_core.vhd:451:33  */
  assign decoder_b_n147 = decoder_b_clk_multi_cycle_o; // (signal)
  /* upi41_core.vhd:452:33  */
  assign decoder_b_n148 = decoder_b_clk_assert_psen_o; // (signal)
  /* upi41_core.vhd:453:33  */
  assign decoder_b_n149 = decoder_b_clk_assert_prog_o; // (signal)
  /* upi41_core.vhd:454:33  */
  assign decoder_b_n150 = decoder_b_clk_assert_rd_o; // (signal)
  /* upi41_core.vhd:455:33  */
  assign decoder_b_n151 = decoder_b_clk_assert_wr_o; // (signal)
  /* upi41_core.vhd:458:33  */
  assign decoder_b_n152 = decoder_b_cnd_compute_take_o; // (signal)
  /* upi41_core.vhd:459:33  */
  assign decoder_b_n153 = decoder_b_cnd_branch_cond_o; // (signal)
  /* upi41_core.vhd:461:33  */
  assign decoder_b_n154 = decoder_b_cnd_comp_value_o; // (signal)
  /* upi41_core.vhd:462:33  */
  assign decoder_b_n155 = decoder_b_cnd_f1_o; // (signal)
  /* upi41_core.vhd:463:33  */
  assign decoder_b_n156 = decoder_b_cnd_tf_o; // (signal)
  /* upi41_core.vhd:464:33  */
  assign decoder_b_n157 = decoder_b_dm_addr_type_o; // (signal)
  /* upi41_core.vhd:465:33  */
  assign decoder_b_n158 = decoder_b_tim_read_timer_o; // (signal)
  /* upi41_core.vhd:466:33  */
  assign decoder_b_n159 = decoder_b_tim_write_timer_o; // (signal)
  /* upi41_core.vhd:467:33  */
  assign decoder_b_n160 = decoder_b_tim_start_t_o; // (signal)
  /* upi41_core.vhd:468:33  */
  assign decoder_b_n161 = decoder_b_tim_start_cnt_o; // (signal)
  /* upi41_core.vhd:469:33  */
  assign decoder_b_n162 = decoder_b_tim_stop_tcnt_o; // (signal)
  /* upi41_core.vhd:470:33  */
  assign decoder_b_n163 = decoder_b_p1_read_reg_o; // (signal)
  /* upi41_core.vhd:471:33  */
  assign decoder_b_n164 = decoder_b_p2_read_reg_o; // (signal)
  /* upi41_core.vhd:472:33  */
  assign decoder_b_n165 = decoder_b_p2_read_exp_o; // (signal)
  /* upi41_core.vhd:473:33  */
  assign decoder_b_n166 = decoder_b_p2_output_pch_o; // (signal)
  /* upi41_core.vhd:474:33  */
  assign decoder_b_n167 = decoder_b_pm_inc_pc_o; // (signal)
  /* upi41_core.vhd:475:33  */
  assign decoder_b_n168 = decoder_b_pm_write_pmem_addr_o; // (signal)
  /* upi41_core.vhd:476:33  */
  assign decoder_b_n169 = decoder_b_pm_addr_type_o; // (signal)
  /* upi41_core.vhd:477:33  */
  assign decoder_b_n170 = decoder_b_psw_special_data_o; // (signal)
  /* upi41_core.vhd:481:33  */
  assign decoder_b_n171 = decoder_b_psw_inc_stackp_o; // (signal)
  /* upi41_core.vhd:482:33  */
  assign decoder_b_n172 = decoder_b_psw_dec_stackp_o; // (signal)
  /* upi41_core.vhd:483:33  */
  assign decoder_b_n173 = decoder_b_psw_write_carry_o; // (signal)
  /* upi41_core.vhd:484:33  */
  assign decoder_b_n174 = decoder_b_psw_write_aux_carry_o; // (signal)
  /* upi41_core.vhd:485:33  */
  assign decoder_b_n175 = decoder_b_psw_write_f0_o; // (signal)
  /* upi41_core.vhd:486:33  */
  assign decoder_b_n176 = decoder_b_psw_write_bs_o; // (signal)
  /* upi41_core.vhd:394:3  */
  t48_decoder_1_1_1 decoder_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_s),
    .ea_i(gnd_s),
    .ale_i(ale_s),
    .int_n_i(bus_int_n_s),
    .data_i(t48_data_s),
    .bus_set_f1_i(bus_set_f1_s),
    .bus_clear_f1_i(bus_clear_f1_s),
    .alu_carry_i(alu_carry_s),
    .alu_da_overflow_i(alu_da_overflow_s),
    .clk_mstate_i(clk_mstate_s),
    .clk_second_cycle_i(clk_second_cycle_s),
    .cnd_take_branch_i(cnd_take_branch_s),
    .psw_carry_i(psw_carry_s),
    .psw_aux_carry_i(psw_aux_carry_s),
    .psw_f0_i(psw_f0_s),
    .tim_overflow_i(tim_overflow_s),
    .t0_dir_o(),
    .data_o(decoder_b_data_o),
    .alu_write_accu_o(decoder_b_alu_write_accu_o),
    .alu_write_shadow_o(decoder_b_alu_write_shadow_o),
    .alu_write_temp_reg_o(decoder_b_alu_write_temp_reg_o),
    .alu_read_alu_o(decoder_b_alu_read_alu_o),
    .bus_write_bus_o(decoder_b_bus_write_bus_o),
    .bus_read_bus_o(decoder_b_bus_read_bus_o),
    .bus_ibf_int_o(decoder_b_bus_ibf_int_o),
    .bus_en_dma_o(decoder_b_bus_en_dma_o),
    .bus_en_flags_o(decoder_b_bus_en_flags_o),
    .bus_write_sts_o(decoder_b_bus_write_sts_o),
    .dm_write_dmem_addr_o(decoder_b_dm_write_dmem_addr_o),
    .dm_write_dmem_o(decoder_b_dm_write_dmem_o),
    .dm_read_dmem_o(decoder_b_dm_read_dmem_o),
    .p1_write_p1_o(decoder_b_p1_write_p1_o),
    .p1_read_p1_o(decoder_b_p1_read_p1_o),
    .p2_write_p2_o(decoder_b_p2_write_p2_o),
    .p2_write_exp_o(decoder_b_p2_write_exp_o),
    .p2_read_p2_o(decoder_b_p2_read_p2_o),
    .p2_read_exp_o(decoder_b_p2_read_exp_o),
    .pm_write_pcl_o(decoder_b_pm_write_pcl_o),
    .pm_read_pcl_o(decoder_b_pm_read_pcl_o),
    .pm_write_pch_o(decoder_b_pm_write_pch_o),
    .pm_read_pch_o(decoder_b_pm_read_pch_o),
    .pm_read_pmem_o(decoder_b_pm_read_pmem_o),
    .psw_read_psw_o(decoder_b_psw_read_psw_o),
    .psw_read_sp_o(decoder_b_psw_read_sp_o),
    .psw_write_psw_o(decoder_b_psw_write_psw_o),
    .psw_write_sp_o(decoder_b_psw_write_sp_o),
    .alu_op_o(decoder_b_alu_op_o),
    .alu_use_carry_o(decoder_b_alu_use_carry_o),
    .alu_da_high_o(decoder_b_alu_da_high_o),
    .alu_accu_low_o(decoder_b_alu_accu_low_o),
    .alu_p06_temp_reg_o(decoder_b_alu_p06_temp_reg_o),
    .alu_p60_temp_reg_o(decoder_b_alu_p60_temp_reg_o),
    .bus_output_pcl_o(),
    .bus_bidir_bus_o(),
    .clk_multi_cycle_o(decoder_b_clk_multi_cycle_o),
    .clk_assert_psen_o(decoder_b_clk_assert_psen_o),
    .clk_assert_prog_o(decoder_b_clk_assert_prog_o),
    .clk_assert_rd_o(decoder_b_clk_assert_rd_o),
    .clk_assert_wr_o(decoder_b_clk_assert_wr_o),
    .cnd_compute_take_o(decoder_b_cnd_compute_take_o),
    .cnd_branch_cond_o(decoder_b_cnd_branch_cond_o),
    .cnd_comp_value_o(decoder_b_cnd_comp_value_o),
    .cnd_f1_o(decoder_b_cnd_f1_o),
    .cnd_tf_o(decoder_b_cnd_tf_o),
    .dm_addr_type_o(decoder_b_dm_addr_type_o),
    .p1_read_reg_o(decoder_b_p1_read_reg_o),
    .p2_read_reg_o(decoder_b_p2_read_reg_o),
    .p2_output_pch_o(decoder_b_p2_output_pch_o),
    .pm_inc_pc_o(decoder_b_pm_inc_pc_o),
    .pm_write_pmem_addr_o(decoder_b_pm_write_pmem_addr_o),
    .pm_addr_type_o(decoder_b_pm_addr_type_o),
    .psw_special_data_o(decoder_b_psw_special_data_o),
    .psw_inc_stackp_o(decoder_b_psw_inc_stackp_o),
    .psw_dec_stackp_o(decoder_b_psw_dec_stackp_o),
    .psw_write_carry_o(decoder_b_psw_write_carry_o),
    .psw_write_aux_carry_o(decoder_b_psw_write_aux_carry_o),
    .psw_write_f0_o(decoder_b_psw_write_f0_o),
    .psw_write_bs_o(decoder_b_psw_write_bs_o),
    .tim_read_timer_o(decoder_b_tim_read_timer_o),
    .tim_write_timer_o(decoder_b_tim_write_timer_o),
    .tim_start_t_o(decoder_b_tim_start_t_o),
    .tim_start_cnt_o(decoder_b_tim_start_cnt_o),
    .tim_stop_tcnt_o(decoder_b_tim_stop_tcnt_o));
  /* upi41_core.vhd:501:28  */
  assign dmem_ctrl_b_n308 = dmem_ctrl_b_data_o; // (signal)
  /* upi41_core.vhd:503:28  */
  assign dmem_ctrl_b_n309 = dmem_ctrl_b_dmem_addr_o; // (signal)
  /* upi41_core.vhd:504:28  */
  assign dmem_ctrl_b_n310 = dmem_ctrl_b_dmem_we_o; // (signal)
  /* upi41_core.vhd:505:28  */
  assign dmem_ctrl_b_n311 = dmem_ctrl_b_dmem_data_o; // (signal)
  /* upi41_core.vhd:490:3  */
  t48_dmem_ctrl dmem_ctrl_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_dmem_addr_i(dm_write_dmem_addr_s),
    .write_dmem_i(dm_write_dmem_s),
    .read_dmem_i(dm_read_dmem_s),
    .addr_type_i(dm_addr_type_s),
    .bank_select_i(psw_bs_s),
    .dmem_data_i(dmem_data_i),
    .data_o(dmem_ctrl_b_data_o),
    .dmem_addr_o(dmem_ctrl_b_dmem_addr_o),
    .dmem_we_o(dmem_ctrl_b_dmem_we_o),
    .dmem_data_o(dmem_ctrl_b_dmem_data_o));
  /* upi41_core.vhd:519:24  */
  assign timer_b_n320 = timer_b_data_o; // (signal)
  /* upi41_core.vhd:525:24  */
  assign timer_b_n321 = timer_b_overflow_o; // (signal)
  /* upi41_core.vhd:508:3  */
  t48_timer_4 timer_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .t1_i(t1_s),
    .clk_mstate_i(clk_mstate_s),
    .data_i(t48_data_s),
    .read_timer_i(tim_read_timer_s),
    .write_timer_i(tim_write_timer_s),
    .start_t_i(tim_start_t_s),
    .start_cnt_i(tim_start_cnt_s),
    .stop_tcnt_i(tim_stop_tcnt_s),
    .data_o(timer_b_data_o),
    .overflow_o(timer_b_overflow_o));
  /* t48_pack-p.vhd:75:5  */
  assign n333_o = tim_of_s ? 1'b1 : 1'b0;
  /* upi41_core.vhd:536:23  */
  assign p1_b_n334 = p1_b_data_o; // (signal)
  /* upi41_core.vhd:541:23  */
  assign p1_b_n335 = p1_b_p1_o; // (signal)
  /* upi41_core.vhd:542:23  */
  assign p1_b_n336 = p1_b_p1_low_imp_o; // (signal)
  /* upi41_core.vhd:530:3  */
  t48_p1 p1_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_p1_i(p1_write_p1_s),
    .read_p1_i(p1_read_p1_s),
    .read_reg_i(p1_read_reg_s),
    .p1_i(p1_i),
    .data_o(p1_b_data_o),
    .p1_o(p1_b_p1_o),
    .p1_low_imp_o(p1_b_p1_low_imp_o));
  /* upi41_core.vhd:553:24  */
  assign p2_b_n343 = p2_b_data_o; // (signal)
  /* upi41_core.vhd:560:35  */
  assign n344_o = pmem_addr_s[11:8];
  /* upi41_core.vhd:562:24  */
  assign p2_b_n345 = p2_b_p2_o; // (signal)
  /* upi41_core.vhd:563:24  */
  assign p2_b_n346 = p2_b_p2l_low_imp_o; // (signal)
  /* upi41_core.vhd:564:24  */
  assign p2_b_n347 = p2_b_p2h_low_imp_o; // (signal)
  /* upi41_core.vhd:545:3  */
  t48_p2 p2_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_s),
    .data_i(t48_data_s),
    .write_p2_i(p2_write_p2_s),
    .write_exp_i(p2_write_exp_s),
    .read_p2_i(p2_read_p2_s),
    .read_reg_i(p2_read_reg_s),
    .read_exp_i(p2_read_exp_s),
    .output_pch_i(p2_output_pch_s),
    .pch_i(n344_o),
    .p2_i(p2_i),
    .data_o(p2_b_data_o),
    .p2_o(p2_b_p2_o),
    .p2l_low_imp_o(p2_b_p2l_low_imp_o),
    .p2h_low_imp_o(p2_b_p2h_low_imp_o));
  /* upi41_core.vhd:567:16  */
  assign n356_o = p2_s[6];
  /* upi41_core.vhd:567:25  */
  assign n357_o = ~bus_dma_s;
  /* upi41_core.vhd:567:20  */
  assign n358_o = n357_o ? n356_o : bus_drq_s;
  /* upi41_core.vhd:568:17  */
  assign n359_o = p2_s[7];
  /* upi41_core.vhd:569:11  */
  assign n360_o = {n359_o, p26_s};
  /* upi41_core.vhd:570:18  */
  assign n361_o = p2_s[5];
  /* upi41_core.vhd:570:22  */
  assign n362_o = n361_o & bus_mint_ibf_n_s;
  /* upi41_core.vhd:570:11  */
  assign n363_o = {n360_o, n362_o};
  /* upi41_core.vhd:571:18  */
  assign n364_o = p2_s[4];
  /* upi41_core.vhd:571:22  */
  assign n365_o = n364_o & bus_mint_obf_s;
  /* upi41_core.vhd:571:11  */
  assign n366_o = {n363_o, n365_o};
  /* upi41_core.vhd:572:17  */
  assign n367_o = p2_s[3:0];
  /* upi41_core.vhd:572:11  */
  assign n368_o = {n366_o, n367_o};
  /* upi41_core.vhd:580:28  */
  assign pmem_ctrl_b_n369 = pmem_ctrl_b_data_o; // (signal)
  /* upi41_core.vhd:589:28  */
  assign pmem_ctrl_b_n370 = pmem_ctrl_b_pmem_addr_o; // (signal)
  /* upi41_core.vhd:574:3  */
  t48_pmem_ctrl pmem_ctrl_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_pcl_i(pm_write_pcl_s),
    .read_pcl_i(pm_read_pcl_s),
    .write_pch_i(pm_write_pch_s),
    .read_pch_i(pm_read_pch_s),
    .inc_pc_i(pm_inc_pc_s),
    .write_pmem_addr_i(pm_write_pmem_addr_s),
    .addr_type_i(pm_addr_type_s),
    .read_pmem_i(pm_read_pmem_s),
    .pmem_data_i(pmem_data_i),
    .data_o(pmem_ctrl_b_data_o),
    .pmem_addr_o(pmem_ctrl_b_pmem_addr_o));
  /* upi41_core.vhd:599:29  */
  assign psw_b_n375 = psw_b_data_o; // (signal)
  /* upi41_core.vhd:611:29  */
  assign psw_b_n376 = psw_b_carry_o; // (signal)
  /* upi41_core.vhd:613:29  */
  assign psw_b_n377 = psw_b_aux_carry_o; // (signal)
  /* upi41_core.vhd:614:29  */
  assign psw_b_n378 = psw_b_f0_o; // (signal)
  /* upi41_core.vhd:615:29  */
  assign psw_b_n379 = psw_b_bs_o; // (signal)
  /* upi41_core.vhd:593:3  */
  t48_psw psw_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .read_psw_i(psw_read_psw_s),
    .read_sp_i(psw_read_sp_s),
    .write_psw_i(psw_write_psw_s),
    .write_sp_i(psw_write_sp_s),
    .special_data_i(psw_special_data_s),
    .inc_stackp_i(psw_inc_stackp_s),
    .dec_stackp_i(psw_dec_stackp_s),
    .write_carry_i(psw_write_carry_s),
    .write_aux_carry_i(psw_write_aux_carry_s),
    .write_f0_i(psw_write_f0_s),
    .write_bs_i(psw_write_bs_s),
    .aux_carry_i(alu_aux_carry_s),
    .data_o(psw_b_data_o),
    .carry_o(psw_b_carry_o),
    .aux_carry_o(psw_b_aux_carry_o),
    .f0_o(psw_b_f0_o),
    .bs_o(psw_b_bs_o));
  /* upi41_core.vhd:622:30  */
  assign n391_o = ~prog_s;
  /* t48_pack-p.vhd:66:5  */
  assign n398_o = n391_o ? 1'b1 : 1'b0;
  /* t48_pack-p.vhd:66:5  */
  assign n406_o = xtal3_s ? 1'b1 : 1'b0;
  /* upi41_core.vhd:624:29  */
  assign n407_o = pmem_addr_s[10:0];
endmodule

