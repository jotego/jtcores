
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"cc",x"fa",x"c2",x"87"),
    12 => (x"86",x"c0",x"c5",x"4e"),
    13 => (x"49",x"cc",x"fa",x"c2"),
    14 => (x"48",x"c0",x"e7",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e7",x"e0"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"71",x"1e",x"4f",x"26"),
    53 => (x"49",x"66",x"c4",x"4a"),
    54 => (x"c8",x"88",x"c1",x"48"),
    55 => (x"99",x"71",x"58",x"a6"),
    56 => (x"ff",x"87",x"d6",x"02"),
    57 => (x"ff",x"c3",x"48",x"d4"),
    58 => (x"c4",x"52",x"68",x"78"),
    59 => (x"c1",x"48",x"49",x"66"),
    60 => (x"58",x"a6",x"c8",x"88"),
    61 => (x"ea",x"05",x"99",x"71"),
    62 => (x"1e",x"4f",x"26",x"87"),
    63 => (x"d4",x"ff",x"1e",x"73"),
    64 => (x"7b",x"ff",x"c3",x"4b"),
    65 => (x"ff",x"c3",x"4a",x"6b"),
    66 => (x"c8",x"49",x"6b",x"7b"),
    67 => (x"c3",x"b1",x"72",x"32"),
    68 => (x"4a",x"6b",x"7b",x"ff"),
    69 => (x"b2",x"71",x"31",x"c8"),
    70 => (x"6b",x"7b",x"ff",x"c3"),
    71 => (x"72",x"32",x"c8",x"49"),
    72 => (x"c4",x"48",x"71",x"b1"),
    73 => (x"26",x"4d",x"26",x"87"),
    74 => (x"26",x"4b",x"26",x"4c"),
    75 => (x"5b",x"5e",x"0e",x"4f"),
    76 => (x"71",x"0e",x"5d",x"5c"),
    77 => (x"4c",x"d4",x"ff",x"4a"),
    78 => (x"ff",x"c3",x"49",x"72"),
    79 => (x"c2",x"7c",x"71",x"99"),
    80 => (x"05",x"bf",x"c0",x"e7"),
    81 => (x"66",x"d0",x"87",x"c8"),
    82 => (x"d4",x"30",x"c9",x"48"),
    83 => (x"66",x"d0",x"58",x"a6"),
    84 => (x"c3",x"29",x"d8",x"49"),
    85 => (x"7c",x"71",x"99",x"ff"),
    86 => (x"d0",x"49",x"66",x"d0"),
    87 => (x"99",x"ff",x"c3",x"29"),
    88 => (x"66",x"d0",x"7c",x"71"),
    89 => (x"c3",x"29",x"c8",x"49"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"c3",x"49",x"66",x"d0"),
    92 => (x"7c",x"71",x"99",x"ff"),
    93 => (x"29",x"d0",x"49",x"72"),
    94 => (x"71",x"99",x"ff",x"c3"),
    95 => (x"c9",x"4b",x"6c",x"7c"),
    96 => (x"c3",x"4d",x"ff",x"f0"),
    97 => (x"d0",x"05",x"ab",x"ff"),
    98 => (x"7c",x"ff",x"c3",x"87"),
    99 => (x"8d",x"c1",x"4b",x"6c"),
   100 => (x"c3",x"87",x"c6",x"02"),
   101 => (x"f0",x"02",x"ab",x"ff"),
   102 => (x"fe",x"48",x"73",x"87"),
   103 => (x"c0",x"1e",x"87",x"c7"),
   104 => (x"48",x"d4",x"ff",x"49"),
   105 => (x"c1",x"78",x"ff",x"c3"),
   106 => (x"b7",x"c8",x"c3",x"81"),
   107 => (x"87",x"f1",x"04",x"a9"),
   108 => (x"73",x"1e",x"4f",x"26"),
   109 => (x"c4",x"87",x"e7",x"1e"),
   110 => (x"c0",x"4b",x"df",x"f8"),
   111 => (x"f0",x"ff",x"c0",x"1e"),
   112 => (x"fd",x"49",x"f7",x"c1"),
   113 => (x"86",x"c4",x"87",x"e7"),
   114 => (x"c0",x"05",x"a8",x"c1"),
   115 => (x"d4",x"ff",x"87",x"ea"),
   116 => (x"78",x"ff",x"c3",x"48"),
   117 => (x"c0",x"c0",x"c0",x"c1"),
   118 => (x"c0",x"1e",x"c0",x"c0"),
   119 => (x"e9",x"c1",x"f0",x"e1"),
   120 => (x"87",x"c9",x"fd",x"49"),
   121 => (x"98",x"70",x"86",x"c4"),
   122 => (x"ff",x"87",x"ca",x"05"),
   123 => (x"ff",x"c3",x"48",x"d4"),
   124 => (x"cb",x"48",x"c1",x"78"),
   125 => (x"87",x"e6",x"fe",x"87"),
   126 => (x"fe",x"05",x"8b",x"c1"),
   127 => (x"48",x"c0",x"87",x"fd"),
   128 => (x"1e",x"87",x"e6",x"fc"),
   129 => (x"d4",x"ff",x"1e",x"73"),
   130 => (x"78",x"ff",x"c3",x"48"),
   131 => (x"1e",x"c0",x"4b",x"d3"),
   132 => (x"c1",x"f0",x"ff",x"c0"),
   133 => (x"d4",x"fc",x"49",x"c1"),
   134 => (x"70",x"86",x"c4",x"87"),
   135 => (x"87",x"ca",x"05",x"98"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"48",x"c1",x"78",x"ff"),
   138 => (x"f1",x"fd",x"87",x"cb"),
   139 => (x"05",x"8b",x"c1",x"87"),
   140 => (x"c0",x"87",x"db",x"ff"),
   141 => (x"87",x"f1",x"fb",x"48"),
   142 => (x"5c",x"5b",x"5e",x"0e"),
   143 => (x"4c",x"d4",x"ff",x"0e"),
   144 => (x"c6",x"87",x"db",x"fd"),
   145 => (x"e1",x"c0",x"1e",x"ea"),
   146 => (x"49",x"c8",x"c1",x"f0"),
   147 => (x"c4",x"87",x"de",x"fb"),
   148 => (x"02",x"a8",x"c1",x"86"),
   149 => (x"ea",x"fe",x"87",x"c8"),
   150 => (x"c1",x"48",x"c0",x"87"),
   151 => (x"da",x"fa",x"87",x"e2"),
   152 => (x"cf",x"49",x"70",x"87"),
   153 => (x"c6",x"99",x"ff",x"ff"),
   154 => (x"c8",x"02",x"a9",x"ea"),
   155 => (x"87",x"d3",x"fe",x"87"),
   156 => (x"cb",x"c1",x"48",x"c0"),
   157 => (x"7c",x"ff",x"c3",x"87"),
   158 => (x"fc",x"4b",x"f1",x"c0"),
   159 => (x"98",x"70",x"87",x"f4"),
   160 => (x"87",x"eb",x"c0",x"02"),
   161 => (x"ff",x"c0",x"1e",x"c0"),
   162 => (x"49",x"fa",x"c1",x"f0"),
   163 => (x"c4",x"87",x"de",x"fa"),
   164 => (x"05",x"98",x"70",x"86"),
   165 => (x"ff",x"c3",x"87",x"d9"),
   166 => (x"c3",x"49",x"6c",x"7c"),
   167 => (x"7c",x"7c",x"7c",x"ff"),
   168 => (x"99",x"c0",x"c1",x"7c"),
   169 => (x"c1",x"87",x"c4",x"02"),
   170 => (x"c0",x"87",x"d5",x"48"),
   171 => (x"c2",x"87",x"d1",x"48"),
   172 => (x"87",x"c4",x"05",x"ab"),
   173 => (x"87",x"c8",x"48",x"c0"),
   174 => (x"fe",x"05",x"8b",x"c1"),
   175 => (x"48",x"c0",x"87",x"fd"),
   176 => (x"1e",x"87",x"e4",x"f9"),
   177 => (x"e7",x"c2",x"1e",x"73"),
   178 => (x"78",x"c1",x"48",x"c0"),
   179 => (x"d0",x"ff",x"4b",x"c7"),
   180 => (x"fb",x"78",x"c2",x"48"),
   181 => (x"d0",x"ff",x"87",x"c8"),
   182 => (x"c0",x"78",x"c3",x"48"),
   183 => (x"d0",x"e5",x"c0",x"1e"),
   184 => (x"f9",x"49",x"c0",x"c1"),
   185 => (x"86",x"c4",x"87",x"c7"),
   186 => (x"c1",x"05",x"a8",x"c1"),
   187 => (x"ab",x"c2",x"4b",x"87"),
   188 => (x"c0",x"87",x"c5",x"05"),
   189 => (x"87",x"f9",x"c0",x"48"),
   190 => (x"ff",x"05",x"8b",x"c1"),
   191 => (x"f7",x"fc",x"87",x"d0"),
   192 => (x"c4",x"e7",x"c2",x"87"),
   193 => (x"05",x"98",x"70",x"58"),
   194 => (x"1e",x"c1",x"87",x"cd"),
   195 => (x"c1",x"f0",x"ff",x"c0"),
   196 => (x"d8",x"f8",x"49",x"d0"),
   197 => (x"ff",x"86",x"c4",x"87"),
   198 => (x"ff",x"c3",x"48",x"d4"),
   199 => (x"87",x"fc",x"c2",x"78"),
   200 => (x"58",x"c8",x"e7",x"c2"),
   201 => (x"c2",x"48",x"d0",x"ff"),
   202 => (x"48",x"d4",x"ff",x"78"),
   203 => (x"c1",x"78",x"ff",x"c3"),
   204 => (x"87",x"f5",x"f7",x"48"),
   205 => (x"5c",x"5b",x"5e",x"0e"),
   206 => (x"4b",x"71",x"0e",x"5d"),
   207 => (x"ee",x"c5",x"4c",x"c0"),
   208 => (x"ff",x"4a",x"df",x"cd"),
   209 => (x"ff",x"c3",x"48",x"d4"),
   210 => (x"c3",x"49",x"68",x"78"),
   211 => (x"c0",x"05",x"a9",x"fe"),
   212 => (x"4d",x"70",x"87",x"fd"),
   213 => (x"cc",x"02",x"9b",x"73"),
   214 => (x"1e",x"66",x"d0",x"87"),
   215 => (x"f1",x"f5",x"49",x"73"),
   216 => (x"d6",x"86",x"c4",x"87"),
   217 => (x"48",x"d0",x"ff",x"87"),
   218 => (x"c3",x"78",x"d1",x"c4"),
   219 => (x"66",x"d0",x"7d",x"ff"),
   220 => (x"d4",x"88",x"c1",x"48"),
   221 => (x"98",x"70",x"58",x"a6"),
   222 => (x"ff",x"87",x"f0",x"05"),
   223 => (x"ff",x"c3",x"48",x"d4"),
   224 => (x"9b",x"73",x"78",x"78"),
   225 => (x"ff",x"87",x"c5",x"05"),
   226 => (x"78",x"d0",x"48",x"d0"),
   227 => (x"c1",x"4c",x"4a",x"c1"),
   228 => (x"ee",x"fe",x"05",x"8a"),
   229 => (x"f6",x"48",x"74",x"87"),
   230 => (x"73",x"1e",x"87",x"cb"),
   231 => (x"c0",x"4a",x"71",x"1e"),
   232 => (x"48",x"d4",x"ff",x"4b"),
   233 => (x"ff",x"78",x"ff",x"c3"),
   234 => (x"c3",x"c4",x"48",x"d0"),
   235 => (x"48",x"d4",x"ff",x"78"),
   236 => (x"72",x"78",x"ff",x"c3"),
   237 => (x"f0",x"ff",x"c0",x"1e"),
   238 => (x"f5",x"49",x"d1",x"c1"),
   239 => (x"86",x"c4",x"87",x"ef"),
   240 => (x"d2",x"05",x"98",x"70"),
   241 => (x"1e",x"c0",x"c8",x"87"),
   242 => (x"fd",x"49",x"66",x"cc"),
   243 => (x"86",x"c4",x"87",x"e6"),
   244 => (x"d0",x"ff",x"4b",x"70"),
   245 => (x"73",x"78",x"c2",x"48"),
   246 => (x"87",x"cd",x"f5",x"48"),
   247 => (x"5c",x"5b",x"5e",x"0e"),
   248 => (x"1e",x"c0",x"0e",x"5d"),
   249 => (x"c1",x"f0",x"ff",x"c0"),
   250 => (x"c0",x"f5",x"49",x"c9"),
   251 => (x"c2",x"1e",x"d2",x"87"),
   252 => (x"fc",x"49",x"c8",x"e7"),
   253 => (x"86",x"c8",x"87",x"fe"),
   254 => (x"84",x"c1",x"4c",x"c0"),
   255 => (x"04",x"ac",x"b7",x"d2"),
   256 => (x"e7",x"c2",x"87",x"f8"),
   257 => (x"49",x"bf",x"97",x"c8"),
   258 => (x"c1",x"99",x"c0",x"c3"),
   259 => (x"c0",x"05",x"a9",x"c0"),
   260 => (x"e7",x"c2",x"87",x"e7"),
   261 => (x"49",x"bf",x"97",x"cf"),
   262 => (x"e7",x"c2",x"31",x"d0"),
   263 => (x"4a",x"bf",x"97",x"d0"),
   264 => (x"b1",x"72",x"32",x"c8"),
   265 => (x"97",x"d1",x"e7",x"c2"),
   266 => (x"71",x"b1",x"4a",x"bf"),
   267 => (x"ff",x"ff",x"cf",x"4c"),
   268 => (x"84",x"c1",x"9c",x"ff"),
   269 => (x"e7",x"c1",x"34",x"ca"),
   270 => (x"d1",x"e7",x"c2",x"87"),
   271 => (x"c1",x"49",x"bf",x"97"),
   272 => (x"c2",x"99",x"c6",x"31"),
   273 => (x"bf",x"97",x"d2",x"e7"),
   274 => (x"2a",x"b7",x"c7",x"4a"),
   275 => (x"e7",x"c2",x"b1",x"72"),
   276 => (x"4a",x"bf",x"97",x"cd"),
   277 => (x"c2",x"9d",x"cf",x"4d"),
   278 => (x"bf",x"97",x"ce",x"e7"),
   279 => (x"ca",x"9a",x"c3",x"4a"),
   280 => (x"cf",x"e7",x"c2",x"32"),
   281 => (x"c2",x"4b",x"bf",x"97"),
   282 => (x"c2",x"b2",x"73",x"33"),
   283 => (x"bf",x"97",x"d0",x"e7"),
   284 => (x"9b",x"c0",x"c3",x"4b"),
   285 => (x"73",x"2b",x"b7",x"c6"),
   286 => (x"c1",x"81",x"c2",x"b2"),
   287 => (x"70",x"30",x"71",x"48"),
   288 => (x"75",x"48",x"c1",x"49"),
   289 => (x"72",x"4d",x"70",x"30"),
   290 => (x"71",x"84",x"c1",x"4c"),
   291 => (x"b7",x"c0",x"c8",x"94"),
   292 => (x"87",x"cc",x"06",x"ad"),
   293 => (x"2d",x"b7",x"34",x"c1"),
   294 => (x"ad",x"b7",x"c0",x"c8"),
   295 => (x"87",x"f4",x"ff",x"01"),
   296 => (x"c0",x"f2",x"48",x"74"),
   297 => (x"5b",x"5e",x"0e",x"87"),
   298 => (x"f8",x"0e",x"5d",x"5c"),
   299 => (x"ee",x"ef",x"c2",x"86"),
   300 => (x"c2",x"78",x"c0",x"48"),
   301 => (x"c0",x"1e",x"e6",x"e7"),
   302 => (x"87",x"de",x"fb",x"49"),
   303 => (x"98",x"70",x"86",x"c4"),
   304 => (x"c0",x"87",x"c5",x"05"),
   305 => (x"87",x"ce",x"c9",x"48"),
   306 => (x"7e",x"c1",x"4d",x"c0"),
   307 => (x"bf",x"da",x"f5",x"c0"),
   308 => (x"dc",x"e8",x"c2",x"49"),
   309 => (x"4b",x"c8",x"71",x"4a"),
   310 => (x"70",x"87",x"cf",x"ee"),
   311 => (x"87",x"c2",x"05",x"98"),
   312 => (x"f5",x"c0",x"7e",x"c0"),
   313 => (x"c2",x"49",x"bf",x"d6"),
   314 => (x"71",x"4a",x"f8",x"e8"),
   315 => (x"f9",x"ed",x"4b",x"c8"),
   316 => (x"05",x"98",x"70",x"87"),
   317 => (x"7e",x"c0",x"87",x"c2"),
   318 => (x"fd",x"c0",x"02",x"6e"),
   319 => (x"ec",x"ee",x"c2",x"87"),
   320 => (x"ef",x"c2",x"4d",x"bf"),
   321 => (x"7e",x"bf",x"9f",x"e4"),
   322 => (x"ea",x"d6",x"c5",x"48"),
   323 => (x"87",x"c7",x"05",x"a8"),
   324 => (x"bf",x"ec",x"ee",x"c2"),
   325 => (x"6e",x"87",x"ce",x"4d"),
   326 => (x"d5",x"e9",x"ca",x"48"),
   327 => (x"87",x"c5",x"02",x"a8"),
   328 => (x"f1",x"c7",x"48",x"c0"),
   329 => (x"e6",x"e7",x"c2",x"87"),
   330 => (x"f9",x"49",x"75",x"1e"),
   331 => (x"86",x"c4",x"87",x"ec"),
   332 => (x"c5",x"05",x"98",x"70"),
   333 => (x"c7",x"48",x"c0",x"87"),
   334 => (x"f5",x"c0",x"87",x"dc"),
   335 => (x"c2",x"49",x"bf",x"d6"),
   336 => (x"71",x"4a",x"f8",x"e8"),
   337 => (x"e1",x"ec",x"4b",x"c8"),
   338 => (x"05",x"98",x"70",x"87"),
   339 => (x"ef",x"c2",x"87",x"c8"),
   340 => (x"78",x"c1",x"48",x"ee"),
   341 => (x"f5",x"c0",x"87",x"da"),
   342 => (x"c2",x"49",x"bf",x"da"),
   343 => (x"71",x"4a",x"dc",x"e8"),
   344 => (x"c5",x"ec",x"4b",x"c8"),
   345 => (x"02",x"98",x"70",x"87"),
   346 => (x"c0",x"87",x"c5",x"c0"),
   347 => (x"87",x"e6",x"c6",x"48"),
   348 => (x"97",x"e4",x"ef",x"c2"),
   349 => (x"d5",x"c1",x"49",x"bf"),
   350 => (x"cd",x"c0",x"05",x"a9"),
   351 => (x"e5",x"ef",x"c2",x"87"),
   352 => (x"c2",x"49",x"bf",x"97"),
   353 => (x"c0",x"02",x"a9",x"ea"),
   354 => (x"48",x"c0",x"87",x"c5"),
   355 => (x"c2",x"87",x"c7",x"c6"),
   356 => (x"bf",x"97",x"e6",x"e7"),
   357 => (x"e9",x"c3",x"48",x"7e"),
   358 => (x"ce",x"c0",x"02",x"a8"),
   359 => (x"c3",x"48",x"6e",x"87"),
   360 => (x"c0",x"02",x"a8",x"eb"),
   361 => (x"48",x"c0",x"87",x"c5"),
   362 => (x"c2",x"87",x"eb",x"c5"),
   363 => (x"bf",x"97",x"f1",x"e7"),
   364 => (x"c0",x"05",x"99",x"49"),
   365 => (x"e7",x"c2",x"87",x"cc"),
   366 => (x"49",x"bf",x"97",x"f2"),
   367 => (x"c0",x"02",x"a9",x"c2"),
   368 => (x"48",x"c0",x"87",x"c5"),
   369 => (x"c2",x"87",x"cf",x"c5"),
   370 => (x"bf",x"97",x"f3",x"e7"),
   371 => (x"ea",x"ef",x"c2",x"48"),
   372 => (x"48",x"4c",x"70",x"58"),
   373 => (x"ef",x"c2",x"88",x"c1"),
   374 => (x"e7",x"c2",x"58",x"ee"),
   375 => (x"49",x"bf",x"97",x"f4"),
   376 => (x"e7",x"c2",x"81",x"75"),
   377 => (x"4a",x"bf",x"97",x"f5"),
   378 => (x"a1",x"72",x"32",x"c8"),
   379 => (x"fb",x"f3",x"c2",x"7e"),
   380 => (x"c2",x"78",x"6e",x"48"),
   381 => (x"bf",x"97",x"f6",x"e7"),
   382 => (x"58",x"a6",x"c8",x"48"),
   383 => (x"bf",x"ee",x"ef",x"c2"),
   384 => (x"87",x"d4",x"c2",x"02"),
   385 => (x"bf",x"d6",x"f5",x"c0"),
   386 => (x"f8",x"e8",x"c2",x"49"),
   387 => (x"4b",x"c8",x"71",x"4a"),
   388 => (x"70",x"87",x"d7",x"e9"),
   389 => (x"c5",x"c0",x"02",x"98"),
   390 => (x"c3",x"48",x"c0",x"87"),
   391 => (x"ef",x"c2",x"87",x"f8"),
   392 => (x"c2",x"4c",x"bf",x"e6"),
   393 => (x"c2",x"5c",x"cf",x"f4"),
   394 => (x"bf",x"97",x"cb",x"e8"),
   395 => (x"c2",x"31",x"c8",x"49"),
   396 => (x"bf",x"97",x"ca",x"e8"),
   397 => (x"c2",x"49",x"a1",x"4a"),
   398 => (x"bf",x"97",x"cc",x"e8"),
   399 => (x"72",x"32",x"d0",x"4a"),
   400 => (x"e8",x"c2",x"49",x"a1"),
   401 => (x"4a",x"bf",x"97",x"cd"),
   402 => (x"a1",x"72",x"32",x"d8"),
   403 => (x"91",x"66",x"c4",x"49"),
   404 => (x"bf",x"fb",x"f3",x"c2"),
   405 => (x"c3",x"f4",x"c2",x"81"),
   406 => (x"d3",x"e8",x"c2",x"59"),
   407 => (x"c8",x"4a",x"bf",x"97"),
   408 => (x"d2",x"e8",x"c2",x"32"),
   409 => (x"a2",x"4b",x"bf",x"97"),
   410 => (x"d4",x"e8",x"c2",x"4a"),
   411 => (x"d0",x"4b",x"bf",x"97"),
   412 => (x"4a",x"a2",x"73",x"33"),
   413 => (x"97",x"d5",x"e8",x"c2"),
   414 => (x"9b",x"cf",x"4b",x"bf"),
   415 => (x"a2",x"73",x"33",x"d8"),
   416 => (x"c7",x"f4",x"c2",x"4a"),
   417 => (x"c3",x"f4",x"c2",x"5a"),
   418 => (x"8a",x"c2",x"4a",x"bf"),
   419 => (x"f4",x"c2",x"92",x"74"),
   420 => (x"a1",x"72",x"48",x"c7"),
   421 => (x"87",x"ca",x"c1",x"78"),
   422 => (x"97",x"f8",x"e7",x"c2"),
   423 => (x"31",x"c8",x"49",x"bf"),
   424 => (x"97",x"f7",x"e7",x"c2"),
   425 => (x"49",x"a1",x"4a",x"bf"),
   426 => (x"59",x"f6",x"ef",x"c2"),
   427 => (x"bf",x"f2",x"ef",x"c2"),
   428 => (x"c7",x"31",x"c5",x"49"),
   429 => (x"29",x"c9",x"81",x"ff"),
   430 => (x"59",x"cf",x"f4",x"c2"),
   431 => (x"97",x"fd",x"e7",x"c2"),
   432 => (x"32",x"c8",x"4a",x"bf"),
   433 => (x"97",x"fc",x"e7",x"c2"),
   434 => (x"4a",x"a2",x"4b",x"bf"),
   435 => (x"6e",x"92",x"66",x"c4"),
   436 => (x"cb",x"f4",x"c2",x"82"),
   437 => (x"c3",x"f4",x"c2",x"5a"),
   438 => (x"c2",x"78",x"c0",x"48"),
   439 => (x"72",x"48",x"ff",x"f3"),
   440 => (x"f4",x"c2",x"78",x"a1"),
   441 => (x"f4",x"c2",x"48",x"cf"),
   442 => (x"c2",x"78",x"bf",x"c3"),
   443 => (x"c2",x"48",x"d3",x"f4"),
   444 => (x"78",x"bf",x"c7",x"f4"),
   445 => (x"bf",x"ee",x"ef",x"c2"),
   446 => (x"87",x"c9",x"c0",x"02"),
   447 => (x"30",x"c4",x"48",x"74"),
   448 => (x"c9",x"c0",x"7e",x"70"),
   449 => (x"cb",x"f4",x"c2",x"87"),
   450 => (x"30",x"c4",x"48",x"bf"),
   451 => (x"ef",x"c2",x"7e",x"70"),
   452 => (x"78",x"6e",x"48",x"f2"),
   453 => (x"8e",x"f8",x"48",x"c1"),
   454 => (x"4c",x"26",x"4d",x"26"),
   455 => (x"4f",x"26",x"4b",x"26"),
   456 => (x"5c",x"5b",x"5e",x"0e"),
   457 => (x"4a",x"71",x"0e",x"5d"),
   458 => (x"bf",x"ee",x"ef",x"c2"),
   459 => (x"72",x"87",x"cb",x"02"),
   460 => (x"72",x"2b",x"c7",x"4b"),
   461 => (x"9c",x"ff",x"c1",x"4c"),
   462 => (x"4b",x"72",x"87",x"c9"),
   463 => (x"4c",x"72",x"2b",x"c8"),
   464 => (x"c2",x"9c",x"ff",x"c3"),
   465 => (x"83",x"bf",x"fb",x"f3"),
   466 => (x"bf",x"d2",x"f5",x"c0"),
   467 => (x"87",x"d9",x"02",x"ab"),
   468 => (x"5b",x"d6",x"f5",x"c0"),
   469 => (x"1e",x"e6",x"e7",x"c2"),
   470 => (x"fd",x"f0",x"49",x"73"),
   471 => (x"70",x"86",x"c4",x"87"),
   472 => (x"87",x"c5",x"05",x"98"),
   473 => (x"e6",x"c0",x"48",x"c0"),
   474 => (x"ee",x"ef",x"c2",x"87"),
   475 => (x"87",x"d2",x"02",x"bf"),
   476 => (x"91",x"c4",x"49",x"74"),
   477 => (x"81",x"e6",x"e7",x"c2"),
   478 => (x"ff",x"cf",x"4d",x"69"),
   479 => (x"9d",x"ff",x"ff",x"ff"),
   480 => (x"49",x"74",x"87",x"cb"),
   481 => (x"e7",x"c2",x"91",x"c2"),
   482 => (x"69",x"9f",x"81",x"e6"),
   483 => (x"fe",x"48",x"75",x"4d"),
   484 => (x"5e",x"0e",x"87",x"c6"),
   485 => (x"0e",x"5d",x"5c",x"5b"),
   486 => (x"c0",x"4d",x"71",x"1e"),
   487 => (x"cf",x"49",x"c1",x"1e"),
   488 => (x"86",x"c4",x"87",x"d4"),
   489 => (x"02",x"9c",x"4c",x"70"),
   490 => (x"c2",x"87",x"c0",x"c1"),
   491 => (x"75",x"4a",x"f6",x"ef"),
   492 => (x"87",x"db",x"e2",x"49"),
   493 => (x"c0",x"02",x"98",x"70"),
   494 => (x"4a",x"74",x"87",x"f1"),
   495 => (x"4b",x"cb",x"49",x"75"),
   496 => (x"70",x"87",x"c1",x"e3"),
   497 => (x"e2",x"c0",x"02",x"98"),
   498 => (x"74",x"1e",x"c0",x"87"),
   499 => (x"87",x"c7",x"02",x"9c"),
   500 => (x"c0",x"48",x"a6",x"c4"),
   501 => (x"c4",x"87",x"c5",x"78"),
   502 => (x"78",x"c1",x"48",x"a6"),
   503 => (x"ce",x"49",x"66",x"c4"),
   504 => (x"86",x"c4",x"87",x"d4"),
   505 => (x"05",x"9c",x"4c",x"70"),
   506 => (x"74",x"87",x"c0",x"ff"),
   507 => (x"e7",x"fc",x"26",x"48"),
   508 => (x"5b",x"5e",x"0e",x"87"),
   509 => (x"1e",x"0e",x"5d",x"5c"),
   510 => (x"05",x"9b",x"4b",x"71"),
   511 => (x"48",x"c0",x"87",x"c5"),
   512 => (x"c8",x"87",x"e5",x"c1"),
   513 => (x"7d",x"c0",x"4d",x"a3"),
   514 => (x"c7",x"02",x"66",x"d4"),
   515 => (x"97",x"66",x"d4",x"87"),
   516 => (x"87",x"c5",x"05",x"bf"),
   517 => (x"cf",x"c1",x"48",x"c0"),
   518 => (x"49",x"66",x"d4",x"87"),
   519 => (x"70",x"87",x"f3",x"fd"),
   520 => (x"c1",x"02",x"9c",x"4c"),
   521 => (x"a4",x"dc",x"87",x"c0"),
   522 => (x"da",x"7d",x"69",x"49"),
   523 => (x"a3",x"c4",x"49",x"a4"),
   524 => (x"7a",x"69",x"9f",x"4a"),
   525 => (x"bf",x"ee",x"ef",x"c2"),
   526 => (x"d4",x"87",x"d2",x"02"),
   527 => (x"69",x"9f",x"49",x"a4"),
   528 => (x"ff",x"ff",x"c0",x"49"),
   529 => (x"d0",x"48",x"71",x"99"),
   530 => (x"c2",x"7e",x"70",x"30"),
   531 => (x"6e",x"7e",x"c0",x"87"),
   532 => (x"80",x"6a",x"48",x"49"),
   533 => (x"7b",x"c0",x"7a",x"70"),
   534 => (x"6a",x"49",x"a3",x"cc"),
   535 => (x"49",x"a3",x"d0",x"79"),
   536 => (x"48",x"74",x"79",x"c0"),
   537 => (x"48",x"c0",x"87",x"c2"),
   538 => (x"87",x"ec",x"fa",x"26"),
   539 => (x"5c",x"5b",x"5e",x"0e"),
   540 => (x"4c",x"71",x"0e",x"5d"),
   541 => (x"ca",x"c1",x"02",x"9c"),
   542 => (x"49",x"a4",x"c8",x"87"),
   543 => (x"c2",x"c1",x"02",x"69"),
   544 => (x"4a",x"66",x"d0",x"87"),
   545 => (x"d4",x"82",x"49",x"6c"),
   546 => (x"66",x"d0",x"5a",x"a6"),
   547 => (x"ef",x"c2",x"b9",x"4d"),
   548 => (x"ff",x"4a",x"bf",x"ea"),
   549 => (x"71",x"99",x"72",x"ba"),
   550 => (x"e4",x"c0",x"02",x"99"),
   551 => (x"4b",x"a4",x"c4",x"87"),
   552 => (x"fb",x"f9",x"49",x"6b"),
   553 => (x"c2",x"7b",x"70",x"87"),
   554 => (x"49",x"bf",x"e6",x"ef"),
   555 => (x"7c",x"71",x"81",x"6c"),
   556 => (x"ef",x"c2",x"b9",x"75"),
   557 => (x"ff",x"4a",x"bf",x"ea"),
   558 => (x"71",x"99",x"72",x"ba"),
   559 => (x"dc",x"ff",x"05",x"99"),
   560 => (x"f9",x"7c",x"75",x"87"),
   561 => (x"73",x"1e",x"87",x"d2"),
   562 => (x"9b",x"4b",x"71",x"1e"),
   563 => (x"c8",x"87",x"c7",x"02"),
   564 => (x"05",x"69",x"49",x"a3"),
   565 => (x"48",x"c0",x"87",x"c5"),
   566 => (x"c2",x"87",x"ef",x"c0"),
   567 => (x"4a",x"bf",x"ff",x"f3"),
   568 => (x"69",x"49",x"a3",x"c4"),
   569 => (x"c2",x"89",x"c2",x"49"),
   570 => (x"91",x"bf",x"e6",x"ef"),
   571 => (x"c2",x"4a",x"a2",x"71"),
   572 => (x"49",x"bf",x"ea",x"ef"),
   573 => (x"a2",x"71",x"99",x"6b"),
   574 => (x"d6",x"f5",x"c0",x"4a"),
   575 => (x"1e",x"66",x"c8",x"5a"),
   576 => (x"d5",x"ea",x"49",x"72"),
   577 => (x"70",x"86",x"c4",x"87"),
   578 => (x"cf",x"f8",x"48",x"49"),
   579 => (x"5b",x"5e",x"0e",x"87"),
   580 => (x"1e",x"0e",x"5d",x"5c"),
   581 => (x"66",x"d4",x"4b",x"71"),
   582 => (x"73",x"2c",x"c9",x"4c"),
   583 => (x"cf",x"c1",x"02",x"9b"),
   584 => (x"49",x"a3",x"c8",x"87"),
   585 => (x"c7",x"c1",x"02",x"69"),
   586 => (x"4d",x"a3",x"d0",x"87"),
   587 => (x"c2",x"7d",x"66",x"d4"),
   588 => (x"49",x"bf",x"ea",x"ef"),
   589 => (x"4a",x"6b",x"b9",x"ff"),
   590 => (x"ac",x"71",x"7e",x"99"),
   591 => (x"c0",x"87",x"cd",x"03"),
   592 => (x"a3",x"cc",x"7d",x"7b"),
   593 => (x"49",x"a3",x"c4",x"4a"),
   594 => (x"87",x"c2",x"79",x"6a"),
   595 => (x"9c",x"74",x"8c",x"72"),
   596 => (x"49",x"87",x"dd",x"02"),
   597 => (x"fc",x"49",x"73",x"1e"),
   598 => (x"86",x"c4",x"87",x"d2"),
   599 => (x"c7",x"49",x"66",x"d4"),
   600 => (x"cb",x"02",x"99",x"ff"),
   601 => (x"e6",x"e7",x"c2",x"87"),
   602 => (x"fd",x"49",x"73",x"1e"),
   603 => (x"86",x"c4",x"87",x"d8"),
   604 => (x"87",x"e4",x"f6",x"26"),
   605 => (x"5c",x"5b",x"5e",x"0e"),
   606 => (x"86",x"f0",x"0e",x"5d"),
   607 => (x"c0",x"59",x"a6",x"d0"),
   608 => (x"cc",x"4b",x"66",x"e4"),
   609 => (x"87",x"ca",x"02",x"66"),
   610 => (x"70",x"80",x"c8",x"48"),
   611 => (x"05",x"bf",x"6e",x"7e"),
   612 => (x"48",x"c0",x"87",x"c5"),
   613 => (x"cc",x"87",x"ec",x"c3"),
   614 => (x"84",x"d0",x"4c",x"66"),
   615 => (x"a6",x"c4",x"49",x"73"),
   616 => (x"c4",x"78",x"6c",x"48"),
   617 => (x"80",x"c4",x"81",x"66"),
   618 => (x"c8",x"78",x"bf",x"6e"),
   619 => (x"c6",x"06",x"a9",x"66"),
   620 => (x"66",x"c4",x"49",x"87"),
   621 => (x"c0",x"4b",x"71",x"89"),
   622 => (x"c4",x"01",x"ab",x"b7"),
   623 => (x"c2",x"c3",x"48",x"87"),
   624 => (x"48",x"66",x"c4",x"87"),
   625 => (x"70",x"98",x"ff",x"c7"),
   626 => (x"c1",x"02",x"6e",x"7e"),
   627 => (x"c0",x"c8",x"87",x"c9"),
   628 => (x"71",x"89",x"6e",x"49"),
   629 => (x"e6",x"e7",x"c2",x"4a"),
   630 => (x"73",x"85",x"6e",x"4d"),
   631 => (x"c1",x"06",x"aa",x"b7"),
   632 => (x"49",x"72",x"4a",x"87"),
   633 => (x"80",x"66",x"c4",x"48"),
   634 => (x"8b",x"72",x"7c",x"70"),
   635 => (x"71",x"8a",x"c1",x"49"),
   636 => (x"87",x"d9",x"02",x"99"),
   637 => (x"48",x"66",x"e0",x"c0"),
   638 => (x"e0",x"c0",x"50",x"15"),
   639 => (x"80",x"c1",x"48",x"66"),
   640 => (x"58",x"a6",x"e4",x"c0"),
   641 => (x"8a",x"c1",x"49",x"72"),
   642 => (x"e7",x"05",x"99",x"71"),
   643 => (x"d0",x"1e",x"c1",x"87"),
   644 => (x"d7",x"f9",x"49",x"66"),
   645 => (x"c0",x"86",x"c4",x"87"),
   646 => (x"c1",x"06",x"ab",x"b7"),
   647 => (x"e0",x"c0",x"87",x"e3"),
   648 => (x"ff",x"c7",x"4d",x"66"),
   649 => (x"c0",x"06",x"ab",x"b7"),
   650 => (x"1e",x"75",x"87",x"e2"),
   651 => (x"fa",x"49",x"66",x"d0"),
   652 => (x"c0",x"c8",x"87",x"d4"),
   653 => (x"c8",x"48",x"6c",x"85"),
   654 => (x"7c",x"70",x"80",x"c0"),
   655 => (x"c1",x"8b",x"c0",x"c8"),
   656 => (x"49",x"66",x"d4",x"1e"),
   657 => (x"c8",x"87",x"e5",x"f8"),
   658 => (x"87",x"ee",x"c0",x"86"),
   659 => (x"1e",x"e6",x"e7",x"c2"),
   660 => (x"f9",x"49",x"66",x"d0"),
   661 => (x"86",x"c4",x"87",x"f0"),
   662 => (x"4a",x"e6",x"e7",x"c2"),
   663 => (x"6c",x"48",x"49",x"73"),
   664 => (x"73",x"7c",x"70",x"80"),
   665 => (x"71",x"8b",x"c1",x"49"),
   666 => (x"87",x"ce",x"02",x"99"),
   667 => (x"c1",x"7d",x"97",x"12"),
   668 => (x"c1",x"49",x"73",x"85"),
   669 => (x"05",x"99",x"71",x"8b"),
   670 => (x"b7",x"c0",x"87",x"f2"),
   671 => (x"e1",x"fe",x"01",x"ab"),
   672 => (x"f0",x"48",x"c1",x"87"),
   673 => (x"87",x"d0",x"f2",x"8e"),
   674 => (x"5c",x"5b",x"5e",x"0e"),
   675 => (x"4b",x"71",x"0e",x"5d"),
   676 => (x"87",x"c7",x"02",x"9b"),
   677 => (x"6d",x"4d",x"a3",x"c8"),
   678 => (x"ff",x"87",x"c5",x"05"),
   679 => (x"87",x"fd",x"c0",x"48"),
   680 => (x"6c",x"4c",x"a3",x"d0"),
   681 => (x"99",x"ff",x"c7",x"49"),
   682 => (x"6c",x"87",x"d8",x"05"),
   683 => (x"c1",x"87",x"c9",x"02"),
   684 => (x"f6",x"49",x"73",x"1e"),
   685 => (x"86",x"c4",x"87",x"f6"),
   686 => (x"1e",x"e6",x"e7",x"c2"),
   687 => (x"c5",x"f8",x"49",x"73"),
   688 => (x"6c",x"86",x"c4",x"87"),
   689 => (x"04",x"aa",x"6d",x"4a"),
   690 => (x"48",x"ff",x"87",x"c4"),
   691 => (x"a2",x"c1",x"87",x"cf"),
   692 => (x"c7",x"49",x"72",x"7c"),
   693 => (x"e7",x"c2",x"99",x"ff"),
   694 => (x"69",x"97",x"81",x"e6"),
   695 => (x"87",x"f8",x"f0",x"48"),
   696 => (x"71",x"1e",x"73",x"1e"),
   697 => (x"c0",x"02",x"9b",x"4b"),
   698 => (x"f4",x"c2",x"87",x"e4"),
   699 => (x"4a",x"73",x"5b",x"d3"),
   700 => (x"ef",x"c2",x"8a",x"c2"),
   701 => (x"92",x"49",x"bf",x"e6"),
   702 => (x"bf",x"ff",x"f3",x"c2"),
   703 => (x"c2",x"80",x"72",x"48"),
   704 => (x"71",x"58",x"d7",x"f4"),
   705 => (x"c2",x"30",x"c4",x"48"),
   706 => (x"c0",x"58",x"f6",x"ef"),
   707 => (x"f4",x"c2",x"87",x"ed"),
   708 => (x"f4",x"c2",x"48",x"cf"),
   709 => (x"c2",x"78",x"bf",x"c3"),
   710 => (x"c2",x"48",x"d3",x"f4"),
   711 => (x"78",x"bf",x"c7",x"f4"),
   712 => (x"bf",x"ee",x"ef",x"c2"),
   713 => (x"c2",x"87",x"c9",x"02"),
   714 => (x"49",x"bf",x"e6",x"ef"),
   715 => (x"87",x"c7",x"31",x"c4"),
   716 => (x"bf",x"cb",x"f4",x"c2"),
   717 => (x"c2",x"31",x"c4",x"49"),
   718 => (x"ef",x"59",x"f6",x"ef"),
   719 => (x"5e",x"0e",x"87",x"de"),
   720 => (x"71",x"0e",x"5c",x"5b"),
   721 => (x"72",x"4b",x"c0",x"4a"),
   722 => (x"e1",x"c0",x"02",x"9a"),
   723 => (x"49",x"a2",x"da",x"87"),
   724 => (x"c2",x"4b",x"69",x"9f"),
   725 => (x"02",x"bf",x"ee",x"ef"),
   726 => (x"a2",x"d4",x"87",x"cf"),
   727 => (x"49",x"69",x"9f",x"49"),
   728 => (x"ff",x"ff",x"c0",x"4c"),
   729 => (x"c2",x"34",x"d0",x"9c"),
   730 => (x"74",x"4c",x"c0",x"87"),
   731 => (x"49",x"73",x"b3",x"49"),
   732 => (x"ee",x"87",x"ed",x"fd"),
   733 => (x"5e",x"0e",x"87",x"e4"),
   734 => (x"0e",x"5d",x"5c",x"5b"),
   735 => (x"4a",x"71",x"86",x"f4"),
   736 => (x"9a",x"72",x"7e",x"c0"),
   737 => (x"c2",x"87",x"d8",x"02"),
   738 => (x"c0",x"48",x"e2",x"e7"),
   739 => (x"da",x"e7",x"c2",x"78"),
   740 => (x"d3",x"f4",x"c2",x"48"),
   741 => (x"e7",x"c2",x"78",x"bf"),
   742 => (x"f4",x"c2",x"48",x"de"),
   743 => (x"c2",x"78",x"bf",x"cf"),
   744 => (x"c0",x"48",x"c3",x"f0"),
   745 => (x"f2",x"ef",x"c2",x"50"),
   746 => (x"e7",x"c2",x"49",x"bf"),
   747 => (x"71",x"4a",x"bf",x"e2"),
   748 => (x"ca",x"c4",x"03",x"aa"),
   749 => (x"cf",x"49",x"72",x"87"),
   750 => (x"ea",x"c0",x"05",x"99"),
   751 => (x"d2",x"f5",x"c0",x"87"),
   752 => (x"da",x"e7",x"c2",x"48"),
   753 => (x"e7",x"c2",x"78",x"bf"),
   754 => (x"e7",x"c2",x"1e",x"e6"),
   755 => (x"c2",x"49",x"bf",x"da"),
   756 => (x"c1",x"48",x"da",x"e7"),
   757 => (x"ff",x"71",x"78",x"a1"),
   758 => (x"c4",x"87",x"ff",x"de"),
   759 => (x"ce",x"f5",x"c0",x"86"),
   760 => (x"e6",x"e7",x"c2",x"48"),
   761 => (x"c0",x"87",x"cc",x"78"),
   762 => (x"48",x"bf",x"ce",x"f5"),
   763 => (x"c0",x"80",x"e0",x"c0"),
   764 => (x"c2",x"58",x"d2",x"f5"),
   765 => (x"48",x"bf",x"e2",x"e7"),
   766 => (x"e7",x"c2",x"80",x"c1"),
   767 => (x"4e",x"27",x"58",x"e6"),
   768 => (x"bf",x"00",x"00",x"0d"),
   769 => (x"9d",x"4d",x"bf",x"97"),
   770 => (x"87",x"e3",x"c2",x"02"),
   771 => (x"02",x"ad",x"e5",x"c3"),
   772 => (x"c0",x"87",x"dc",x"c2"),
   773 => (x"4b",x"bf",x"ce",x"f5"),
   774 => (x"11",x"49",x"a3",x"cb"),
   775 => (x"05",x"ac",x"cf",x"4c"),
   776 => (x"75",x"87",x"d2",x"c1"),
   777 => (x"c1",x"99",x"df",x"49"),
   778 => (x"c2",x"91",x"cd",x"89"),
   779 => (x"c1",x"81",x"f6",x"ef"),
   780 => (x"51",x"12",x"4a",x"a3"),
   781 => (x"12",x"4a",x"a3",x"c3"),
   782 => (x"4a",x"a3",x"c5",x"51"),
   783 => (x"a3",x"c7",x"51",x"12"),
   784 => (x"c9",x"51",x"12",x"4a"),
   785 => (x"51",x"12",x"4a",x"a3"),
   786 => (x"12",x"4a",x"a3",x"ce"),
   787 => (x"4a",x"a3",x"d0",x"51"),
   788 => (x"a3",x"d2",x"51",x"12"),
   789 => (x"d4",x"51",x"12",x"4a"),
   790 => (x"51",x"12",x"4a",x"a3"),
   791 => (x"12",x"4a",x"a3",x"d6"),
   792 => (x"4a",x"a3",x"d8",x"51"),
   793 => (x"a3",x"dc",x"51",x"12"),
   794 => (x"de",x"51",x"12",x"4a"),
   795 => (x"51",x"12",x"4a",x"a3"),
   796 => (x"fa",x"c0",x"7e",x"c1"),
   797 => (x"c8",x"49",x"74",x"87"),
   798 => (x"eb",x"c0",x"05",x"99"),
   799 => (x"d0",x"49",x"74",x"87"),
   800 => (x"87",x"d1",x"05",x"99"),
   801 => (x"c0",x"02",x"66",x"dc"),
   802 => (x"49",x"73",x"87",x"cb"),
   803 => (x"70",x"0f",x"66",x"dc"),
   804 => (x"d3",x"c0",x"02",x"98"),
   805 => (x"c0",x"05",x"6e",x"87"),
   806 => (x"ef",x"c2",x"87",x"c6"),
   807 => (x"50",x"c0",x"48",x"f6"),
   808 => (x"bf",x"ce",x"f5",x"c0"),
   809 => (x"87",x"e1",x"c2",x"48"),
   810 => (x"48",x"c3",x"f0",x"c2"),
   811 => (x"c2",x"7e",x"50",x"c0"),
   812 => (x"49",x"bf",x"f2",x"ef"),
   813 => (x"bf",x"e2",x"e7",x"c2"),
   814 => (x"04",x"aa",x"71",x"4a"),
   815 => (x"c2",x"87",x"f6",x"fb"),
   816 => (x"05",x"bf",x"d3",x"f4"),
   817 => (x"c2",x"87",x"c8",x"c0"),
   818 => (x"02",x"bf",x"ee",x"ef"),
   819 => (x"c2",x"87",x"f8",x"c1"),
   820 => (x"49",x"bf",x"de",x"e7"),
   821 => (x"70",x"87",x"c9",x"e9"),
   822 => (x"e2",x"e7",x"c2",x"49"),
   823 => (x"48",x"a6",x"c4",x"59"),
   824 => (x"bf",x"de",x"e7",x"c2"),
   825 => (x"ee",x"ef",x"c2",x"78"),
   826 => (x"d8",x"c0",x"02",x"bf"),
   827 => (x"49",x"66",x"c4",x"87"),
   828 => (x"ff",x"ff",x"ff",x"cf"),
   829 => (x"02",x"a9",x"99",x"f8"),
   830 => (x"c0",x"87",x"c5",x"c0"),
   831 => (x"87",x"e1",x"c0",x"4c"),
   832 => (x"dc",x"c0",x"4c",x"c1"),
   833 => (x"49",x"66",x"c4",x"87"),
   834 => (x"99",x"f8",x"ff",x"cf"),
   835 => (x"c8",x"c0",x"02",x"a9"),
   836 => (x"48",x"a6",x"c8",x"87"),
   837 => (x"c5",x"c0",x"78",x"c0"),
   838 => (x"48",x"a6",x"c8",x"87"),
   839 => (x"66",x"c8",x"78",x"c1"),
   840 => (x"05",x"9c",x"74",x"4c"),
   841 => (x"c4",x"87",x"e0",x"c0"),
   842 => (x"89",x"c2",x"49",x"66"),
   843 => (x"bf",x"e6",x"ef",x"c2"),
   844 => (x"f3",x"c2",x"91",x"4a"),
   845 => (x"c2",x"4a",x"bf",x"ff"),
   846 => (x"72",x"48",x"da",x"e7"),
   847 => (x"e7",x"c2",x"78",x"a1"),
   848 => (x"78",x"c0",x"48",x"e2"),
   849 => (x"c0",x"87",x"de",x"f9"),
   850 => (x"e7",x"8e",x"f4",x"48"),
   851 => (x"00",x"00",x"87",x"ca"),
   852 => (x"ff",x"ff",x"00",x"00"),
   853 => (x"0d",x"5e",x"ff",x"ff"),
   854 => (x"0d",x"67",x"00",x"00"),
   855 => (x"41",x"46",x"00",x"00"),
   856 => (x"20",x"32",x"33",x"54"),
   857 => (x"46",x"00",x"20",x"20"),
   858 => (x"36",x"31",x"54",x"41"),
   859 => (x"00",x"20",x"20",x"20"),
   860 => (x"d8",x"f4",x"c2",x"1e"),
   861 => (x"a8",x"dd",x"48",x"bf"),
   862 => (x"c0",x"87",x"c9",x"05"),
   863 => (x"70",x"87",x"db",x"fd"),
   864 => (x"87",x"c8",x"4a",x"49"),
   865 => (x"c3",x"48",x"d4",x"ff"),
   866 => (x"4a",x"68",x"78",x"ff"),
   867 => (x"4f",x"26",x"48",x"72"),
   868 => (x"d8",x"f4",x"c2",x"1e"),
   869 => (x"a8",x"dd",x"48",x"bf"),
   870 => (x"c0",x"87",x"c6",x"05"),
   871 => (x"d9",x"87",x"e7",x"fc"),
   872 => (x"48",x"d4",x"ff",x"87"),
   873 => (x"ff",x"78",x"ff",x"c3"),
   874 => (x"e1",x"c8",x"48",x"d0"),
   875 => (x"48",x"d4",x"ff",x"78"),
   876 => (x"f4",x"c2",x"78",x"d4"),
   877 => (x"d4",x"ff",x"48",x"d7"),
   878 => (x"4f",x"26",x"50",x"bf"),
   879 => (x"48",x"d0",x"ff",x"1e"),
   880 => (x"26",x"78",x"e0",x"c0"),
   881 => (x"e7",x"fe",x"1e",x"4f"),
   882 => (x"99",x"49",x"70",x"87"),
   883 => (x"c0",x"87",x"c6",x"02"),
   884 => (x"f1",x"05",x"a9",x"fb"),
   885 => (x"26",x"48",x"71",x"87"),
   886 => (x"5b",x"5e",x"0e",x"4f"),
   887 => (x"4b",x"71",x"0e",x"5c"),
   888 => (x"cb",x"fe",x"4c",x"c0"),
   889 => (x"99",x"49",x"70",x"87"),
   890 => (x"87",x"f9",x"c0",x"02"),
   891 => (x"02",x"a9",x"ec",x"c0"),
   892 => (x"c0",x"87",x"f2",x"c0"),
   893 => (x"c0",x"02",x"a9",x"fb"),
   894 => (x"66",x"cc",x"87",x"eb"),
   895 => (x"c7",x"03",x"ac",x"b7"),
   896 => (x"02",x"66",x"d0",x"87"),
   897 => (x"53",x"71",x"87",x"c2"),
   898 => (x"c2",x"02",x"99",x"71"),
   899 => (x"fd",x"84",x"c1",x"87"),
   900 => (x"49",x"70",x"87",x"de"),
   901 => (x"87",x"cd",x"02",x"99"),
   902 => (x"02",x"a9",x"ec",x"c0"),
   903 => (x"fb",x"c0",x"87",x"c7"),
   904 => (x"d5",x"ff",x"05",x"a9"),
   905 => (x"02",x"66",x"d0",x"87"),
   906 => (x"97",x"c0",x"87",x"c3"),
   907 => (x"a9",x"ec",x"c0",x"7b"),
   908 => (x"74",x"87",x"c4",x"05"),
   909 => (x"74",x"87",x"c5",x"4a"),
   910 => (x"8a",x"0a",x"c0",x"4a"),
   911 => (x"87",x"c2",x"48",x"72"),
   912 => (x"4c",x"26",x"4d",x"26"),
   913 => (x"4f",x"26",x"4b",x"26"),
   914 => (x"87",x"e4",x"fc",x"1e"),
   915 => (x"f0",x"c0",x"49",x"70"),
   916 => (x"ca",x"04",x"a9",x"b7"),
   917 => (x"b7",x"f9",x"c0",x"87"),
   918 => (x"87",x"c3",x"01",x"a9"),
   919 => (x"c1",x"89",x"f0",x"c0"),
   920 => (x"04",x"a9",x"b7",x"c1"),
   921 => (x"da",x"c1",x"87",x"ca"),
   922 => (x"c3",x"01",x"a9",x"b7"),
   923 => (x"89",x"f7",x"c0",x"87"),
   924 => (x"4f",x"26",x"48",x"71"),
   925 => (x"5c",x"5b",x"5e",x"0e"),
   926 => (x"fc",x"4c",x"71",x"0e"),
   927 => (x"1e",x"c1",x"87",x"d2"),
   928 => (x"74",x"1e",x"66",x"d0"),
   929 => (x"87",x"d1",x"fd",x"49"),
   930 => (x"4b",x"70",x"86",x"c8"),
   931 => (x"c0",x"87",x"ed",x"fc"),
   932 => (x"c2",x"03",x"ab",x"b7"),
   933 => (x"cc",x"8b",x"0b",x"87"),
   934 => (x"03",x"ab",x"b7",x"66"),
   935 => (x"a3",x"74",x"87",x"cf"),
   936 => (x"c0",x"83",x"c1",x"49"),
   937 => (x"66",x"cc",x"51",x"e0"),
   938 => (x"f1",x"04",x"ab",x"b7"),
   939 => (x"49",x"a3",x"74",x"87"),
   940 => (x"cd",x"fe",x"51",x"c0"),
   941 => (x"5b",x"5e",x"0e",x"87"),
   942 => (x"4a",x"71",x"0e",x"5c"),
   943 => (x"72",x"4c",x"d4",x"ff"),
   944 => (x"87",x"ea",x"c0",x"49"),
   945 => (x"02",x"9b",x"4b",x"70"),
   946 => (x"8b",x"c1",x"87",x"c2"),
   947 => (x"c8",x"48",x"d0",x"ff"),
   948 => (x"d5",x"c1",x"78",x"c5"),
   949 => (x"c6",x"49",x"73",x"7c"),
   950 => (x"cf",x"e1",x"c2",x"31"),
   951 => (x"48",x"4a",x"bf",x"97"),
   952 => (x"7c",x"70",x"b0",x"71"),
   953 => (x"c4",x"48",x"d0",x"ff"),
   954 => (x"fd",x"48",x"73",x"78"),
   955 => (x"5e",x"0e",x"87",x"d4"),
   956 => (x"0e",x"5d",x"5c",x"5b"),
   957 => (x"4c",x"71",x"86",x"f4"),
   958 => (x"c0",x"48",x"a6",x"c4"),
   959 => (x"7e",x"a4",x"c8",x"78"),
   960 => (x"49",x"bf",x"97",x"6e"),
   961 => (x"05",x"a9",x"c1",x"c1"),
   962 => (x"a4",x"c9",x"87",x"dd"),
   963 => (x"49",x"69",x"97",x"49"),
   964 => (x"05",x"a9",x"d2",x"c1"),
   965 => (x"a4",x"ca",x"87",x"d1"),
   966 => (x"49",x"69",x"97",x"49"),
   967 => (x"05",x"a9",x"c3",x"c1"),
   968 => (x"48",x"df",x"87",x"c5"),
   969 => (x"f9",x"87",x"e1",x"c2"),
   970 => (x"4b",x"c0",x"87",x"e6"),
   971 => (x"97",x"cd",x"ff",x"c0"),
   972 => (x"a9",x"c0",x"49",x"bf"),
   973 => (x"fa",x"87",x"cf",x"04"),
   974 => (x"83",x"c1",x"87",x"cb"),
   975 => (x"97",x"cd",x"ff",x"c0"),
   976 => (x"06",x"ab",x"49",x"bf"),
   977 => (x"ff",x"c0",x"87",x"f1"),
   978 => (x"02",x"bf",x"97",x"cd"),
   979 => (x"df",x"f8",x"87",x"cf"),
   980 => (x"99",x"49",x"70",x"87"),
   981 => (x"c0",x"87",x"c6",x"02"),
   982 => (x"f1",x"05",x"a9",x"ec"),
   983 => (x"f8",x"4b",x"c0",x"87"),
   984 => (x"4d",x"70",x"87",x"ce"),
   985 => (x"cc",x"87",x"c9",x"f8"),
   986 => (x"c3",x"f8",x"58",x"a6"),
   987 => (x"c1",x"4a",x"70",x"87"),
   988 => (x"bf",x"97",x"6e",x"83"),
   989 => (x"c7",x"02",x"ad",x"49"),
   990 => (x"ad",x"ff",x"c0",x"87"),
   991 => (x"87",x"ea",x"c0",x"05"),
   992 => (x"97",x"49",x"a4",x"c9"),
   993 => (x"66",x"c8",x"49",x"69"),
   994 => (x"87",x"c7",x"02",x"a9"),
   995 => (x"a8",x"ff",x"c0",x"48"),
   996 => (x"ca",x"87",x"d7",x"05"),
   997 => (x"69",x"97",x"49",x"a4"),
   998 => (x"c6",x"02",x"aa",x"49"),
   999 => (x"aa",x"ff",x"c0",x"87"),
  1000 => (x"c4",x"87",x"c7",x"05"),
  1001 => (x"78",x"c1",x"48",x"a6"),
  1002 => (x"ec",x"c0",x"87",x"d3"),
  1003 => (x"87",x"c6",x"02",x"ad"),
  1004 => (x"05",x"ad",x"fb",x"c0"),
  1005 => (x"4b",x"c0",x"87",x"c7"),
  1006 => (x"c1",x"48",x"a6",x"c4"),
  1007 => (x"02",x"66",x"c4",x"78"),
  1008 => (x"f7",x"87",x"dc",x"fe"),
  1009 => (x"48",x"73",x"87",x"f6"),
  1010 => (x"f3",x"f9",x"8e",x"f4"),
  1011 => (x"5e",x"0e",x"00",x"87"),
  1012 => (x"0e",x"5d",x"5c",x"5b"),
  1013 => (x"c0",x"4b",x"71",x"1e"),
  1014 => (x"04",x"ab",x"4d",x"4c"),
  1015 => (x"c0",x"87",x"e8",x"c0"),
  1016 => (x"75",x"1e",x"ee",x"fb"),
  1017 => (x"87",x"c4",x"02",x"9d"),
  1018 => (x"87",x"c2",x"4a",x"c0"),
  1019 => (x"49",x"72",x"4a",x"c1"),
  1020 => (x"c4",x"87",x"c3",x"ee"),
  1021 => (x"c1",x"7e",x"70",x"86"),
  1022 => (x"c2",x"05",x"6e",x"84"),
  1023 => (x"c1",x"4c",x"73",x"87"),
  1024 => (x"06",x"ac",x"73",x"85"),
  1025 => (x"6e",x"87",x"d8",x"ff"),
  1026 => (x"4d",x"26",x"26",x"48"),
  1027 => (x"4b",x"26",x"4c",x"26"),
  1028 => (x"5e",x"0e",x"4f",x"26"),
  1029 => (x"0e",x"5d",x"5c",x"5b"),
  1030 => (x"49",x"4c",x"71",x"1e"),
  1031 => (x"f4",x"c2",x"91",x"de"),
  1032 => (x"85",x"71",x"4d",x"f1"),
  1033 => (x"c1",x"02",x"6d",x"97"),
  1034 => (x"f4",x"c2",x"87",x"dd"),
  1035 => (x"74",x"4a",x"bf",x"dc"),
  1036 => (x"fe",x"49",x"72",x"82"),
  1037 => (x"7e",x"70",x"87",x"d8"),
  1038 => (x"f3",x"c0",x"02",x"6e"),
  1039 => (x"e4",x"f4",x"c2",x"87"),
  1040 => (x"cb",x"4a",x"6e",x"4b"),
  1041 => (x"df",x"c1",x"ff",x"49"),
  1042 => (x"cb",x"4b",x"74",x"87"),
  1043 => (x"d8",x"e2",x"c1",x"93"),
  1044 => (x"c1",x"83",x"c4",x"83"),
  1045 => (x"74",x"7b",x"cb",x"c2"),
  1046 => (x"c8",x"cb",x"c1",x"49"),
  1047 => (x"c2",x"7b",x"75",x"87"),
  1048 => (x"bf",x"97",x"f0",x"f4"),
  1049 => (x"f4",x"c2",x"1e",x"49"),
  1050 => (x"df",x"c1",x"49",x"e4"),
  1051 => (x"86",x"c4",x"87",x"d2"),
  1052 => (x"ca",x"c1",x"49",x"74"),
  1053 => (x"49",x"c0",x"87",x"ef"),
  1054 => (x"87",x"ce",x"cc",x"c1"),
  1055 => (x"48",x"d8",x"f4",x"c2"),
  1056 => (x"49",x"c1",x"78",x"c0"),
  1057 => (x"26",x"87",x"c3",x"dd"),
  1058 => (x"4c",x"87",x"ff",x"fd"),
  1059 => (x"69",x"64",x"61",x"6f"),
  1060 => (x"2e",x"2e",x"67",x"6e"),
  1061 => (x"5e",x"0e",x"00",x"2e"),
  1062 => (x"71",x"0e",x"5c",x"5b"),
  1063 => (x"f4",x"c2",x"4a",x"4b"),
  1064 => (x"72",x"82",x"bf",x"dc"),
  1065 => (x"87",x"e6",x"fc",x"49"),
  1066 => (x"02",x"9c",x"4c",x"70"),
  1067 => (x"ea",x"49",x"87",x"c4"),
  1068 => (x"f4",x"c2",x"87",x"cc"),
  1069 => (x"78",x"c0",x"48",x"dc"),
  1070 => (x"cd",x"dc",x"49",x"c1"),
  1071 => (x"87",x"cc",x"fd",x"87"),
  1072 => (x"5c",x"5b",x"5e",x"0e"),
  1073 => (x"86",x"f4",x"0e",x"5d"),
  1074 => (x"4d",x"e6",x"e7",x"c2"),
  1075 => (x"a6",x"c4",x"4c",x"c0"),
  1076 => (x"c2",x"78",x"c0",x"48"),
  1077 => (x"49",x"bf",x"dc",x"f4"),
  1078 => (x"c1",x"06",x"a9",x"c0"),
  1079 => (x"e7",x"c2",x"87",x"c1"),
  1080 => (x"02",x"98",x"48",x"e6"),
  1081 => (x"c0",x"87",x"f8",x"c0"),
  1082 => (x"c8",x"1e",x"ee",x"fb"),
  1083 => (x"87",x"c7",x"02",x"66"),
  1084 => (x"c0",x"48",x"a6",x"c4"),
  1085 => (x"c4",x"87",x"c5",x"78"),
  1086 => (x"78",x"c1",x"48",x"a6"),
  1087 => (x"e9",x"49",x"66",x"c4"),
  1088 => (x"86",x"c4",x"87",x"f4"),
  1089 => (x"84",x"c1",x"4d",x"70"),
  1090 => (x"c1",x"48",x"66",x"c4"),
  1091 => (x"58",x"a6",x"c8",x"80"),
  1092 => (x"bf",x"dc",x"f4",x"c2"),
  1093 => (x"c6",x"03",x"ac",x"49"),
  1094 => (x"05",x"9d",x"75",x"87"),
  1095 => (x"c0",x"87",x"c8",x"ff"),
  1096 => (x"02",x"9d",x"75",x"4c"),
  1097 => (x"c0",x"87",x"e0",x"c3"),
  1098 => (x"c8",x"1e",x"ee",x"fb"),
  1099 => (x"87",x"c7",x"02",x"66"),
  1100 => (x"c0",x"48",x"a6",x"cc"),
  1101 => (x"cc",x"87",x"c5",x"78"),
  1102 => (x"78",x"c1",x"48",x"a6"),
  1103 => (x"e8",x"49",x"66",x"cc"),
  1104 => (x"86",x"c4",x"87",x"f4"),
  1105 => (x"02",x"6e",x"7e",x"70"),
  1106 => (x"6e",x"87",x"e9",x"c2"),
  1107 => (x"97",x"81",x"cb",x"49"),
  1108 => (x"99",x"d0",x"49",x"69"),
  1109 => (x"87",x"d6",x"c1",x"02"),
  1110 => (x"4a",x"d6",x"c2",x"c1"),
  1111 => (x"91",x"cb",x"49",x"74"),
  1112 => (x"81",x"d8",x"e2",x"c1"),
  1113 => (x"81",x"c8",x"79",x"72"),
  1114 => (x"74",x"51",x"ff",x"c3"),
  1115 => (x"c2",x"91",x"de",x"49"),
  1116 => (x"71",x"4d",x"f1",x"f4"),
  1117 => (x"97",x"c1",x"c2",x"85"),
  1118 => (x"49",x"a5",x"c1",x"7d"),
  1119 => (x"c2",x"51",x"e0",x"c0"),
  1120 => (x"bf",x"97",x"f6",x"ef"),
  1121 => (x"c1",x"87",x"d2",x"02"),
  1122 => (x"4b",x"a5",x"c2",x"84"),
  1123 => (x"4a",x"f6",x"ef",x"c2"),
  1124 => (x"fc",x"fe",x"49",x"db"),
  1125 => (x"db",x"c1",x"87",x"d2"),
  1126 => (x"49",x"a5",x"cd",x"87"),
  1127 => (x"84",x"c1",x"51",x"c0"),
  1128 => (x"6e",x"4b",x"a5",x"c2"),
  1129 => (x"fe",x"49",x"cb",x"4a"),
  1130 => (x"c1",x"87",x"fd",x"fb"),
  1131 => (x"c0",x"c1",x"87",x"c6"),
  1132 => (x"49",x"74",x"4a",x"d2"),
  1133 => (x"e2",x"c1",x"91",x"cb"),
  1134 => (x"79",x"72",x"81",x"d8"),
  1135 => (x"97",x"f6",x"ef",x"c2"),
  1136 => (x"87",x"d8",x"02",x"bf"),
  1137 => (x"91",x"de",x"49",x"74"),
  1138 => (x"f4",x"c2",x"84",x"c1"),
  1139 => (x"83",x"71",x"4b",x"f1"),
  1140 => (x"4a",x"f6",x"ef",x"c2"),
  1141 => (x"fb",x"fe",x"49",x"dd"),
  1142 => (x"87",x"d8",x"87",x"ce"),
  1143 => (x"93",x"de",x"4b",x"74"),
  1144 => (x"83",x"f1",x"f4",x"c2"),
  1145 => (x"c0",x"49",x"a3",x"cb"),
  1146 => (x"73",x"84",x"c1",x"51"),
  1147 => (x"49",x"cb",x"4a",x"6e"),
  1148 => (x"87",x"f4",x"fa",x"fe"),
  1149 => (x"c1",x"48",x"66",x"c4"),
  1150 => (x"58",x"a6",x"c8",x"80"),
  1151 => (x"c0",x"03",x"ac",x"c7"),
  1152 => (x"05",x"6e",x"87",x"c5"),
  1153 => (x"74",x"87",x"e0",x"fc"),
  1154 => (x"f7",x"8e",x"f4",x"48"),
  1155 => (x"73",x"1e",x"87",x"fc"),
  1156 => (x"49",x"4b",x"71",x"1e"),
  1157 => (x"e2",x"c1",x"91",x"cb"),
  1158 => (x"a1",x"c8",x"81",x"d8"),
  1159 => (x"cf",x"e1",x"c2",x"4a"),
  1160 => (x"c9",x"50",x"12",x"48"),
  1161 => (x"ff",x"c0",x"4a",x"a1"),
  1162 => (x"50",x"12",x"48",x"cd"),
  1163 => (x"f4",x"c2",x"81",x"ca"),
  1164 => (x"50",x"11",x"48",x"f0"),
  1165 => (x"97",x"f0",x"f4",x"c2"),
  1166 => (x"c0",x"1e",x"49",x"bf"),
  1167 => (x"ff",x"d7",x"c1",x"49"),
  1168 => (x"d8",x"f4",x"c2",x"87"),
  1169 => (x"c1",x"78",x"de",x"48"),
  1170 => (x"87",x"fe",x"d5",x"49"),
  1171 => (x"87",x"fe",x"f6",x"26"),
  1172 => (x"49",x"4a",x"71",x"1e"),
  1173 => (x"e2",x"c1",x"91",x"cb"),
  1174 => (x"81",x"c8",x"81",x"d8"),
  1175 => (x"f4",x"c2",x"48",x"11"),
  1176 => (x"f4",x"c2",x"58",x"dc"),
  1177 => (x"78",x"c0",x"48",x"dc"),
  1178 => (x"dd",x"d5",x"49",x"c1"),
  1179 => (x"1e",x"4f",x"26",x"87"),
  1180 => (x"c4",x"c1",x"49",x"c0"),
  1181 => (x"4f",x"26",x"87",x"d4"),
  1182 => (x"02",x"99",x"71",x"1e"),
  1183 => (x"e3",x"c1",x"87",x"d2"),
  1184 => (x"50",x"c0",x"48",x"ed"),
  1185 => (x"c9",x"c1",x"80",x"f7"),
  1186 => (x"e2",x"c1",x"40",x"d0"),
  1187 => (x"87",x"ce",x"78",x"d1"),
  1188 => (x"48",x"e9",x"e3",x"c1"),
  1189 => (x"78",x"ca",x"e2",x"c1"),
  1190 => (x"c9",x"c1",x"80",x"fc"),
  1191 => (x"4f",x"26",x"78",x"ef"),
  1192 => (x"5c",x"5b",x"5e",x"0e"),
  1193 => (x"4a",x"4c",x"71",x"0e"),
  1194 => (x"e2",x"c1",x"92",x"cb"),
  1195 => (x"a2",x"c8",x"82",x"d8"),
  1196 => (x"4b",x"a2",x"c9",x"49"),
  1197 => (x"1e",x"4b",x"6b",x"97"),
  1198 => (x"1e",x"49",x"69",x"97"),
  1199 => (x"49",x"12",x"82",x"ca"),
  1200 => (x"87",x"f5",x"e4",x"c0"),
  1201 => (x"c1",x"d4",x"49",x"c0"),
  1202 => (x"c1",x"49",x"74",x"87"),
  1203 => (x"f8",x"87",x"d6",x"c1"),
  1204 => (x"87",x"f8",x"f4",x"8e"),
  1205 => (x"71",x"1e",x"73",x"1e"),
  1206 => (x"c3",x"ff",x"49",x"4b"),
  1207 => (x"fe",x"49",x"73",x"87"),
  1208 => (x"e9",x"f4",x"87",x"fe"),
  1209 => (x"1e",x"73",x"1e",x"87"),
  1210 => (x"a3",x"c6",x"4b",x"71"),
  1211 => (x"87",x"db",x"02",x"4a"),
  1212 => (x"d6",x"02",x"8a",x"c1"),
  1213 => (x"c1",x"02",x"8a",x"87"),
  1214 => (x"02",x"8a",x"87",x"da"),
  1215 => (x"8a",x"87",x"fc",x"c0"),
  1216 => (x"87",x"e1",x"c0",x"02"),
  1217 => (x"87",x"cb",x"02",x"8a"),
  1218 => (x"c7",x"87",x"db",x"c1"),
  1219 => (x"87",x"c0",x"fd",x"49"),
  1220 => (x"c2",x"87",x"de",x"c1"),
  1221 => (x"02",x"bf",x"dc",x"f4"),
  1222 => (x"48",x"87",x"cb",x"c1"),
  1223 => (x"f4",x"c2",x"88",x"c1"),
  1224 => (x"c1",x"c1",x"58",x"e0"),
  1225 => (x"e0",x"f4",x"c2",x"87"),
  1226 => (x"f9",x"c0",x"02",x"bf"),
  1227 => (x"dc",x"f4",x"c2",x"87"),
  1228 => (x"80",x"c1",x"48",x"bf"),
  1229 => (x"58",x"e0",x"f4",x"c2"),
  1230 => (x"c2",x"87",x"eb",x"c0"),
  1231 => (x"49",x"bf",x"dc",x"f4"),
  1232 => (x"f4",x"c2",x"89",x"c6"),
  1233 => (x"b7",x"c0",x"59",x"e0"),
  1234 => (x"87",x"da",x"03",x"a9"),
  1235 => (x"48",x"dc",x"f4",x"c2"),
  1236 => (x"87",x"d2",x"78",x"c0"),
  1237 => (x"bf",x"e0",x"f4",x"c2"),
  1238 => (x"c2",x"87",x"cb",x"02"),
  1239 => (x"48",x"bf",x"dc",x"f4"),
  1240 => (x"f4",x"c2",x"80",x"c6"),
  1241 => (x"49",x"c0",x"58",x"e0"),
  1242 => (x"73",x"87",x"df",x"d1"),
  1243 => (x"f4",x"fe",x"c0",x"49"),
  1244 => (x"87",x"da",x"f2",x"87"),
  1245 => (x"71",x"1e",x"73",x"1e"),
  1246 => (x"d8",x"f4",x"c2",x"4b"),
  1247 => (x"c0",x"78",x"dd",x"48"),
  1248 => (x"87",x"c6",x"d1",x"49"),
  1249 => (x"fe",x"c0",x"49",x"73"),
  1250 => (x"c1",x"f2",x"87",x"db"),
  1251 => (x"5b",x"5e",x"0e",x"87"),
  1252 => (x"4c",x"71",x"0e",x"5c"),
  1253 => (x"74",x"1e",x"66",x"cc"),
  1254 => (x"c1",x"93",x"cb",x"4b"),
  1255 => (x"c4",x"83",x"d8",x"e2"),
  1256 => (x"49",x"6a",x"4a",x"a3"),
  1257 => (x"87",x"d0",x"f4",x"fe"),
  1258 => (x"7b",x"ce",x"c8",x"c1"),
  1259 => (x"d4",x"49",x"a3",x"c8"),
  1260 => (x"a3",x"c9",x"51",x"66"),
  1261 => (x"51",x"66",x"d8",x"49"),
  1262 => (x"dc",x"49",x"a3",x"ca"),
  1263 => (x"f1",x"26",x"51",x"66"),
  1264 => (x"5e",x"0e",x"87",x"ca"),
  1265 => (x"0e",x"5d",x"5c",x"5b"),
  1266 => (x"dc",x"86",x"cc",x"ff"),
  1267 => (x"a6",x"c8",x"59",x"a6"),
  1268 => (x"c4",x"78",x"c0",x"48"),
  1269 => (x"66",x"c8",x"c1",x"80"),
  1270 => (x"c1",x"80",x"c4",x"78"),
  1271 => (x"c1",x"80",x"c4",x"78"),
  1272 => (x"e0",x"f4",x"c2",x"78"),
  1273 => (x"c2",x"78",x"c1",x"48"),
  1274 => (x"48",x"bf",x"d8",x"f4"),
  1275 => (x"cb",x"05",x"a8",x"de"),
  1276 => (x"87",x"cc",x"f3",x"87"),
  1277 => (x"a6",x"cc",x"49",x"70"),
  1278 => (x"87",x"ca",x"ce",x"59"),
  1279 => (x"e7",x"87",x"d1",x"e6"),
  1280 => (x"eb",x"e5",x"87",x"c3"),
  1281 => (x"c0",x"4c",x"70",x"87"),
  1282 => (x"c1",x"02",x"ac",x"fb"),
  1283 => (x"66",x"d8",x"87",x"d8"),
  1284 => (x"87",x"ca",x"c1",x"05"),
  1285 => (x"c1",x"1e",x"1e",x"c0"),
  1286 => (x"fb",x"e3",x"c1",x"1e"),
  1287 => (x"fd",x"49",x"c0",x"1e"),
  1288 => (x"86",x"d0",x"87",x"eb"),
  1289 => (x"02",x"ac",x"fb",x"c0"),
  1290 => (x"c4",x"c1",x"87",x"d9"),
  1291 => (x"82",x"c4",x"4a",x"66"),
  1292 => (x"81",x"c7",x"49",x"6a"),
  1293 => (x"1e",x"c1",x"51",x"74"),
  1294 => (x"49",x"6a",x"1e",x"d8"),
  1295 => (x"d8",x"e6",x"81",x"c8"),
  1296 => (x"c1",x"86",x"c8",x"87"),
  1297 => (x"c0",x"48",x"66",x"c8"),
  1298 => (x"87",x"c7",x"01",x"a8"),
  1299 => (x"c1",x"48",x"a6",x"c8"),
  1300 => (x"c1",x"87",x"ce",x"78"),
  1301 => (x"c1",x"48",x"66",x"c8"),
  1302 => (x"58",x"a6",x"d0",x"88"),
  1303 => (x"e4",x"e5",x"87",x"c3"),
  1304 => (x"48",x"a6",x"d0",x"87"),
  1305 => (x"9c",x"74",x"78",x"c2"),
  1306 => (x"87",x"d6",x"cc",x"02"),
  1307 => (x"c1",x"48",x"66",x"c8"),
  1308 => (x"03",x"a8",x"66",x"cc"),
  1309 => (x"c4",x"87",x"cb",x"cc"),
  1310 => (x"78",x"c0",x"48",x"a6"),
  1311 => (x"78",x"c0",x"80",x"d8"),
  1312 => (x"70",x"87",x"ed",x"e3"),
  1313 => (x"48",x"66",x"d8",x"4c"),
  1314 => (x"c6",x"05",x"a8",x"dd"),
  1315 => (x"48",x"a6",x"dc",x"87"),
  1316 => (x"c1",x"78",x"66",x"d8"),
  1317 => (x"c0",x"05",x"ac",x"d0"),
  1318 => (x"d3",x"e3",x"87",x"e8"),
  1319 => (x"87",x"d0",x"e3",x"87"),
  1320 => (x"ec",x"c0",x"4c",x"70"),
  1321 => (x"87",x"c5",x"05",x"ac"),
  1322 => (x"70",x"87",x"da",x"e4"),
  1323 => (x"ac",x"d0",x"c1",x"4c"),
  1324 => (x"d4",x"87",x"c8",x"05"),
  1325 => (x"80",x"c1",x"48",x"66"),
  1326 => (x"c1",x"58",x"a6",x"d8"),
  1327 => (x"ff",x"02",x"ac",x"d0"),
  1328 => (x"e0",x"c0",x"87",x"d8"),
  1329 => (x"66",x"d8",x"48",x"a6"),
  1330 => (x"48",x"66",x"dc",x"78"),
  1331 => (x"a8",x"66",x"e0",x"c0"),
  1332 => (x"87",x"c0",x"ca",x"05"),
  1333 => (x"48",x"a6",x"e4",x"c0"),
  1334 => (x"80",x"c4",x"78",x"c0"),
  1335 => (x"4d",x"74",x"78",x"c0"),
  1336 => (x"02",x"8d",x"fb",x"c0"),
  1337 => (x"c9",x"87",x"c6",x"c9"),
  1338 => (x"87",x"db",x"02",x"8d"),
  1339 => (x"c1",x"02",x"8d",x"c2"),
  1340 => (x"8d",x"c9",x"87",x"f4"),
  1341 => (x"87",x"cb",x"c4",x"02"),
  1342 => (x"c1",x"02",x"8d",x"c4"),
  1343 => (x"8d",x"c1",x"87",x"c1"),
  1344 => (x"87",x"ff",x"c3",x"02"),
  1345 => (x"c8",x"87",x"e0",x"c8"),
  1346 => (x"91",x"cb",x"49",x"66"),
  1347 => (x"81",x"66",x"c4",x"c1"),
  1348 => (x"6a",x"4a",x"a1",x"c4"),
  1349 => (x"c1",x"1e",x"71",x"7e"),
  1350 => (x"c4",x"48",x"fd",x"de"),
  1351 => (x"a1",x"cc",x"49",x"66"),
  1352 => (x"71",x"41",x"20",x"4a"),
  1353 => (x"f8",x"ff",x"05",x"aa"),
  1354 => (x"26",x"51",x"10",x"87"),
  1355 => (x"f4",x"cd",x"c1",x"49"),
  1356 => (x"87",x"d1",x"e2",x"79"),
  1357 => (x"e8",x"c0",x"4c",x"70"),
  1358 => (x"78",x"c1",x"48",x"a6"),
  1359 => (x"c4",x"87",x"ee",x"c7"),
  1360 => (x"f0",x"c0",x"48",x"a6"),
  1361 => (x"87",x"e8",x"e0",x"78"),
  1362 => (x"ec",x"c0",x"4c",x"70"),
  1363 => (x"c3",x"c0",x"02",x"ac"),
  1364 => (x"5c",x"a6",x"c8",x"87"),
  1365 => (x"02",x"ac",x"ec",x"c0"),
  1366 => (x"d3",x"e0",x"87",x"cc"),
  1367 => (x"c0",x"4c",x"70",x"87"),
  1368 => (x"ff",x"05",x"ac",x"ec"),
  1369 => (x"ec",x"c0",x"87",x"f4"),
  1370 => (x"c3",x"c0",x"02",x"ac"),
  1371 => (x"87",x"c0",x"e0",x"87"),
  1372 => (x"d8",x"1e",x"66",x"c4"),
  1373 => (x"d8",x"1e",x"49",x"66"),
  1374 => (x"c1",x"1e",x"49",x"66"),
  1375 => (x"d8",x"1e",x"fb",x"e3"),
  1376 => (x"c8",x"f8",x"49",x"66"),
  1377 => (x"ca",x"1e",x"c0",x"87"),
  1378 => (x"66",x"e0",x"c0",x"1e"),
  1379 => (x"c1",x"91",x"cb",x"49"),
  1380 => (x"d8",x"81",x"66",x"dc"),
  1381 => (x"a1",x"c4",x"48",x"a6"),
  1382 => (x"bf",x"66",x"d8",x"78"),
  1383 => (x"87",x"f9",x"e0",x"49"),
  1384 => (x"b7",x"c0",x"86",x"d8"),
  1385 => (x"ca",x"c1",x"06",x"a8"),
  1386 => (x"de",x"1e",x"c1",x"87"),
  1387 => (x"bf",x"66",x"c8",x"1e"),
  1388 => (x"87",x"e5",x"e0",x"49"),
  1389 => (x"49",x"70",x"86",x"c8"),
  1390 => (x"88",x"08",x"c0",x"48"),
  1391 => (x"58",x"a6",x"ec",x"c0"),
  1392 => (x"06",x"a8",x"b7",x"c0"),
  1393 => (x"c0",x"87",x"ec",x"c0"),
  1394 => (x"dd",x"48",x"66",x"e8"),
  1395 => (x"c0",x"03",x"a8",x"b7"),
  1396 => (x"bf",x"6e",x"87",x"e1"),
  1397 => (x"66",x"e8",x"c0",x"49"),
  1398 => (x"51",x"e0",x"c0",x"81"),
  1399 => (x"49",x"66",x"e8",x"c0"),
  1400 => (x"bf",x"6e",x"81",x"c1"),
  1401 => (x"51",x"c1",x"c2",x"81"),
  1402 => (x"49",x"66",x"e8",x"c0"),
  1403 => (x"bf",x"6e",x"81",x"c2"),
  1404 => (x"d0",x"51",x"c0",x"81"),
  1405 => (x"80",x"c1",x"48",x"66"),
  1406 => (x"48",x"58",x"a6",x"d4"),
  1407 => (x"78",x"c1",x"80",x"d8"),
  1408 => (x"e1",x"87",x"ea",x"c4"),
  1409 => (x"ec",x"c0",x"87",x"c2"),
  1410 => (x"fb",x"e0",x"58",x"a6"),
  1411 => (x"a6",x"f0",x"c0",x"87"),
  1412 => (x"a8",x"ec",x"c0",x"58"),
  1413 => (x"87",x"c9",x"c0",x"05"),
  1414 => (x"e8",x"c0",x"48",x"a6"),
  1415 => (x"c4",x"c0",x"78",x"66"),
  1416 => (x"cb",x"dd",x"ff",x"87"),
  1417 => (x"49",x"66",x"c8",x"87"),
  1418 => (x"c4",x"c1",x"91",x"cb"),
  1419 => (x"80",x"71",x"48",x"66"),
  1420 => (x"c4",x"58",x"a6",x"c8"),
  1421 => (x"82",x"c8",x"4a",x"66"),
  1422 => (x"ca",x"49",x"66",x"c4"),
  1423 => (x"66",x"e8",x"c0",x"81"),
  1424 => (x"66",x"ec",x"c0",x"51"),
  1425 => (x"c0",x"81",x"c1",x"49"),
  1426 => (x"c1",x"89",x"66",x"e8"),
  1427 => (x"70",x"30",x"71",x"48"),
  1428 => (x"71",x"89",x"c1",x"49"),
  1429 => (x"f8",x"c2",x"7a",x"97"),
  1430 => (x"c0",x"49",x"bf",x"cd"),
  1431 => (x"97",x"29",x"66",x"e8"),
  1432 => (x"71",x"48",x"4a",x"6a"),
  1433 => (x"a6",x"f4",x"c0",x"98"),
  1434 => (x"49",x"66",x"c4",x"58"),
  1435 => (x"7e",x"69",x"81",x"c4"),
  1436 => (x"48",x"66",x"e0",x"c0"),
  1437 => (x"02",x"a8",x"66",x"dc"),
  1438 => (x"dc",x"87",x"c8",x"c0"),
  1439 => (x"78",x"c0",x"48",x"a6"),
  1440 => (x"dc",x"87",x"c5",x"c0"),
  1441 => (x"78",x"c1",x"48",x"a6"),
  1442 => (x"c0",x"1e",x"66",x"dc"),
  1443 => (x"66",x"c8",x"1e",x"e0"),
  1444 => (x"c4",x"dd",x"ff",x"49"),
  1445 => (x"70",x"86",x"c8",x"87"),
  1446 => (x"ac",x"b7",x"c0",x"4c"),
  1447 => (x"87",x"d6",x"c1",x"06"),
  1448 => (x"80",x"74",x"48",x"6e"),
  1449 => (x"e0",x"c0",x"7e",x"70"),
  1450 => (x"6e",x"89",x"74",x"49"),
  1451 => (x"fa",x"de",x"c1",x"4b"),
  1452 => (x"e7",x"fe",x"71",x"4a"),
  1453 => (x"48",x"6e",x"87",x"f2"),
  1454 => (x"7e",x"70",x"80",x"c2"),
  1455 => (x"48",x"66",x"e4",x"c0"),
  1456 => (x"e8",x"c0",x"80",x"c1"),
  1457 => (x"f0",x"c0",x"58",x"a6"),
  1458 => (x"81",x"c1",x"49",x"66"),
  1459 => (x"c0",x"02",x"a9",x"70"),
  1460 => (x"4d",x"c0",x"87",x"c5"),
  1461 => (x"c1",x"87",x"c2",x"c0"),
  1462 => (x"c2",x"1e",x"75",x"4d"),
  1463 => (x"e0",x"c0",x"49",x"a4"),
  1464 => (x"70",x"88",x"71",x"48"),
  1465 => (x"66",x"c8",x"1e",x"49"),
  1466 => (x"ec",x"db",x"ff",x"49"),
  1467 => (x"c0",x"86",x"c8",x"87"),
  1468 => (x"ff",x"01",x"a8",x"b7"),
  1469 => (x"e4",x"c0",x"87",x"c6"),
  1470 => (x"d3",x"c0",x"02",x"66"),
  1471 => (x"49",x"66",x"c4",x"87"),
  1472 => (x"e4",x"c0",x"81",x"c9"),
  1473 => (x"66",x"c4",x"51",x"66"),
  1474 => (x"e0",x"ca",x"c1",x"48"),
  1475 => (x"87",x"ce",x"c0",x"78"),
  1476 => (x"c9",x"49",x"66",x"c4"),
  1477 => (x"c4",x"51",x"c2",x"81"),
  1478 => (x"cb",x"c1",x"48",x"66"),
  1479 => (x"e8",x"c0",x"78",x"d4"),
  1480 => (x"78",x"c1",x"48",x"a6"),
  1481 => (x"ff",x"87",x"c6",x"c0"),
  1482 => (x"70",x"87",x"da",x"da"),
  1483 => (x"66",x"e8",x"c0",x"4c"),
  1484 => (x"87",x"f5",x"c0",x"02"),
  1485 => (x"cc",x"48",x"66",x"c8"),
  1486 => (x"c0",x"04",x"a8",x"66"),
  1487 => (x"66",x"c8",x"87",x"cb"),
  1488 => (x"cc",x"80",x"c1",x"48"),
  1489 => (x"e0",x"c0",x"58",x"a6"),
  1490 => (x"48",x"66",x"cc",x"87"),
  1491 => (x"a6",x"d0",x"88",x"c1"),
  1492 => (x"87",x"d5",x"c0",x"58"),
  1493 => (x"05",x"ac",x"c6",x"c1"),
  1494 => (x"d0",x"87",x"c8",x"c0"),
  1495 => (x"80",x"c1",x"48",x"66"),
  1496 => (x"ff",x"58",x"a6",x"d4"),
  1497 => (x"70",x"87",x"de",x"d9"),
  1498 => (x"48",x"66",x"d4",x"4c"),
  1499 => (x"a6",x"d8",x"80",x"c1"),
  1500 => (x"02",x"9c",x"74",x"58"),
  1501 => (x"c8",x"87",x"cb",x"c0"),
  1502 => (x"cc",x"c1",x"48",x"66"),
  1503 => (x"f3",x"04",x"a8",x"66"),
  1504 => (x"d8",x"ff",x"87",x"f5"),
  1505 => (x"66",x"c8",x"87",x"f6"),
  1506 => (x"03",x"a8",x"c7",x"48"),
  1507 => (x"c2",x"87",x"e5",x"c0"),
  1508 => (x"c0",x"48",x"e0",x"f4"),
  1509 => (x"49",x"66",x"c8",x"78"),
  1510 => (x"c4",x"c1",x"91",x"cb"),
  1511 => (x"a1",x"c4",x"81",x"66"),
  1512 => (x"c0",x"4a",x"6a",x"4a"),
  1513 => (x"66",x"c8",x"79",x"52"),
  1514 => (x"cc",x"80",x"c1",x"48"),
  1515 => (x"a8",x"c7",x"58",x"a6"),
  1516 => (x"87",x"db",x"ff",x"04"),
  1517 => (x"e1",x"8e",x"cc",x"ff"),
  1518 => (x"20",x"3a",x"87",x"d0"),
  1519 => (x"50",x"49",x"44",x"00"),
  1520 => (x"69",x"77",x"53",x"20"),
  1521 => (x"65",x"68",x"63",x"74"),
  1522 => (x"73",x"1e",x"00",x"73"),
  1523 => (x"9b",x"4b",x"71",x"1e"),
  1524 => (x"c2",x"87",x"c6",x"02"),
  1525 => (x"c0",x"48",x"dc",x"f4"),
  1526 => (x"c2",x"1e",x"c7",x"78"),
  1527 => (x"49",x"bf",x"dc",x"f4"),
  1528 => (x"d8",x"e2",x"c1",x"1e"),
  1529 => (x"d8",x"f4",x"c2",x"1e"),
  1530 => (x"d5",x"ef",x"49",x"bf"),
  1531 => (x"c2",x"86",x"cc",x"87"),
  1532 => (x"49",x"bf",x"d8",x"f4"),
  1533 => (x"73",x"87",x"c1",x"ea"),
  1534 => (x"87",x"c8",x"02",x"9b"),
  1535 => (x"49",x"d8",x"e2",x"c1"),
  1536 => (x"87",x"f3",x"ed",x"c0"),
  1537 => (x"1e",x"87",x"c7",x"e0"),
  1538 => (x"c1",x"87",x"cf",x"c7"),
  1539 => (x"87",x"fa",x"fe",x"49"),
  1540 => (x"87",x"ef",x"ea",x"fe"),
  1541 => (x"cd",x"02",x"98",x"70"),
  1542 => (x"c8",x"f2",x"fe",x"87"),
  1543 => (x"02",x"98",x"70",x"87"),
  1544 => (x"4a",x"c1",x"87",x"c4"),
  1545 => (x"4a",x"c0",x"87",x"c2"),
  1546 => (x"ce",x"05",x"9a",x"72"),
  1547 => (x"c1",x"1e",x"c0",x"87"),
  1548 => (x"c0",x"49",x"dc",x"e1"),
  1549 => (x"c4",x"87",x"de",x"f9"),
  1550 => (x"c1",x"87",x"fe",x"86"),
  1551 => (x"c0",x"87",x"fa",x"c0"),
  1552 => (x"e7",x"e1",x"c1",x"1e"),
  1553 => (x"cc",x"f9",x"c0",x"49"),
  1554 => (x"c1",x"1e",x"c0",x"87"),
  1555 => (x"70",x"87",x"c0",x"c3"),
  1556 => (x"c0",x"f9",x"c0",x"49"),
  1557 => (x"87",x"c1",x"c3",x"87"),
  1558 => (x"4f",x"26",x"8e",x"f8"),
  1559 => (x"66",x"20",x"44",x"53"),
  1560 => (x"65",x"6c",x"69",x"61"),
  1561 => (x"42",x"00",x"2e",x"64"),
  1562 => (x"69",x"74",x"6f",x"6f"),
  1563 => (x"2e",x"2e",x"67",x"6e"),
  1564 => (x"c2",x"1e",x"00",x"2e"),
  1565 => (x"c0",x"48",x"dc",x"f4"),
  1566 => (x"d8",x"f4",x"c2",x"78"),
  1567 => (x"fe",x"78",x"c0",x"48"),
  1568 => (x"c4",x"c1",x"87",x"c5"),
  1569 => (x"48",x"c0",x"87",x"e6"),
  1570 => (x"20",x"80",x"4f",x"26"),
  1571 => (x"74",x"69",x"78",x"45"),
  1572 => (x"42",x"20",x"80",x"00"),
  1573 => (x"00",x"6b",x"63",x"61"),
  1574 => (x"00",x"00",x"12",x"50"),
  1575 => (x"00",x"00",x"2d",x"31"),
  1576 => (x"50",x"00",x"00",x"00"),
  1577 => (x"4f",x"00",x"00",x"12"),
  1578 => (x"00",x"00",x"00",x"2d"),
  1579 => (x"12",x"50",x"00",x"00"),
  1580 => (x"2d",x"6d",x"00",x"00"),
  1581 => (x"00",x"00",x"00",x"00"),
  1582 => (x"00",x"12",x"50",x"00"),
  1583 => (x"00",x"2d",x"8b",x"00"),
  1584 => (x"00",x"00",x"00",x"00"),
  1585 => (x"00",x"00",x"12",x"50"),
  1586 => (x"00",x"00",x"2d",x"a9"),
  1587 => (x"50",x"00",x"00",x"00"),
  1588 => (x"c7",x"00",x"00",x"12"),
  1589 => (x"00",x"00",x"00",x"2d"),
  1590 => (x"12",x"50",x"00",x"00"),
  1591 => (x"2d",x"e5",x"00",x"00"),
  1592 => (x"00",x"00",x"00",x"00"),
  1593 => (x"00",x"12",x"50",x"00"),
  1594 => (x"00",x"00",x"00",x"00"),
  1595 => (x"00",x"00",x"00",x"00"),
  1596 => (x"00",x"00",x"12",x"e5"),
  1597 => (x"00",x"00",x"00",x"00"),
  1598 => (x"4c",x"00",x"00",x"00"),
  1599 => (x"20",x"64",x"61",x"6f"),
  1600 => (x"1e",x"00",x"2e",x"2a"),
  1601 => (x"c0",x"48",x"f0",x"fe"),
  1602 => (x"79",x"09",x"cd",x"78"),
  1603 => (x"1e",x"4f",x"26",x"09"),
  1604 => (x"bf",x"f0",x"fe",x"1e"),
  1605 => (x"26",x"26",x"48",x"7e"),
  1606 => (x"f0",x"fe",x"1e",x"4f"),
  1607 => (x"26",x"78",x"c1",x"48"),
  1608 => (x"f0",x"fe",x"1e",x"4f"),
  1609 => (x"26",x"78",x"c0",x"48"),
  1610 => (x"4a",x"71",x"1e",x"4f"),
  1611 => (x"26",x"52",x"52",x"c0"),
  1612 => (x"5b",x"5e",x"0e",x"4f"),
  1613 => (x"f4",x"0e",x"5d",x"5c"),
  1614 => (x"97",x"4d",x"71",x"86"),
  1615 => (x"a5",x"c1",x"7e",x"6d"),
  1616 => (x"48",x"6c",x"97",x"4c"),
  1617 => (x"6e",x"58",x"a6",x"c8"),
  1618 => (x"a8",x"66",x"c4",x"48"),
  1619 => (x"ff",x"87",x"c5",x"05"),
  1620 => (x"87",x"e6",x"c0",x"48"),
  1621 => (x"c2",x"87",x"ca",x"ff"),
  1622 => (x"6c",x"97",x"49",x"a5"),
  1623 => (x"4b",x"a3",x"71",x"4b"),
  1624 => (x"97",x"4b",x"6b",x"97"),
  1625 => (x"48",x"6e",x"7e",x"6c"),
  1626 => (x"a6",x"c8",x"80",x"c1"),
  1627 => (x"cc",x"98",x"c7",x"58"),
  1628 => (x"97",x"70",x"58",x"a6"),
  1629 => (x"87",x"e1",x"fe",x"7c"),
  1630 => (x"8e",x"f4",x"48",x"73"),
  1631 => (x"4c",x"26",x"4d",x"26"),
  1632 => (x"4f",x"26",x"4b",x"26"),
  1633 => (x"5c",x"5b",x"5e",x"0e"),
  1634 => (x"71",x"86",x"f4",x"0e"),
  1635 => (x"4a",x"66",x"d8",x"4c"),
  1636 => (x"c2",x"9a",x"ff",x"c3"),
  1637 => (x"6c",x"97",x"4b",x"a4"),
  1638 => (x"49",x"a1",x"73",x"49"),
  1639 => (x"6c",x"97",x"51",x"72"),
  1640 => (x"c1",x"48",x"6e",x"7e"),
  1641 => (x"58",x"a6",x"c8",x"80"),
  1642 => (x"a6",x"cc",x"98",x"c7"),
  1643 => (x"f4",x"54",x"70",x"58"),
  1644 => (x"87",x"ca",x"ff",x"8e"),
  1645 => (x"e8",x"fd",x"1e",x"1e"),
  1646 => (x"4a",x"bf",x"e0",x"87"),
  1647 => (x"c0",x"e0",x"c0",x"49"),
  1648 => (x"87",x"cb",x"02",x"99"),
  1649 => (x"f8",x"c2",x"1e",x"72"),
  1650 => (x"f7",x"fe",x"49",x"c3"),
  1651 => (x"fc",x"86",x"c4",x"87"),
  1652 => (x"7e",x"70",x"87",x"fd"),
  1653 => (x"26",x"87",x"c2",x"fd"),
  1654 => (x"c2",x"1e",x"4f",x"26"),
  1655 => (x"fd",x"49",x"c3",x"f8"),
  1656 => (x"e6",x"c1",x"87",x"c7"),
  1657 => (x"da",x"fc",x"49",x"f4"),
  1658 => (x"87",x"c8",x"c4",x"87"),
  1659 => (x"ff",x"1e",x"4f",x"26"),
  1660 => (x"e1",x"c8",x"48",x"d0"),
  1661 => (x"48",x"d4",x"ff",x"78"),
  1662 => (x"66",x"c4",x"78",x"c5"),
  1663 => (x"c3",x"87",x"c3",x"02"),
  1664 => (x"66",x"c8",x"78",x"e0"),
  1665 => (x"ff",x"87",x"c6",x"02"),
  1666 => (x"f0",x"c3",x"48",x"d4"),
  1667 => (x"48",x"d4",x"ff",x"78"),
  1668 => (x"d0",x"ff",x"78",x"71"),
  1669 => (x"78",x"e1",x"c8",x"48"),
  1670 => (x"26",x"78",x"e0",x"c0"),
  1671 => (x"5b",x"5e",x"0e",x"4f"),
  1672 => (x"4c",x"71",x"0e",x"5c"),
  1673 => (x"49",x"c3",x"f8",x"c2"),
  1674 => (x"70",x"87",x"c6",x"fc"),
  1675 => (x"aa",x"b7",x"c0",x"4a"),
  1676 => (x"87",x"e3",x"c2",x"04"),
  1677 => (x"05",x"aa",x"e0",x"c3"),
  1678 => (x"eb",x"c1",x"87",x"c9"),
  1679 => (x"78",x"c1",x"48",x"e7"),
  1680 => (x"c3",x"87",x"d4",x"c2"),
  1681 => (x"c9",x"05",x"aa",x"f0"),
  1682 => (x"e3",x"eb",x"c1",x"87"),
  1683 => (x"c1",x"78",x"c1",x"48"),
  1684 => (x"eb",x"c1",x"87",x"f5"),
  1685 => (x"c7",x"02",x"bf",x"e7"),
  1686 => (x"c2",x"4b",x"72",x"87"),
  1687 => (x"87",x"c2",x"b3",x"c0"),
  1688 => (x"9c",x"74",x"4b",x"72"),
  1689 => (x"c1",x"87",x"d1",x"05"),
  1690 => (x"1e",x"bf",x"e3",x"eb"),
  1691 => (x"bf",x"e7",x"eb",x"c1"),
  1692 => (x"fd",x"49",x"72",x"1e"),
  1693 => (x"86",x"c8",x"87",x"f8"),
  1694 => (x"bf",x"e3",x"eb",x"c1"),
  1695 => (x"87",x"e0",x"c0",x"02"),
  1696 => (x"b7",x"c4",x"49",x"73"),
  1697 => (x"ed",x"c1",x"91",x"29"),
  1698 => (x"4a",x"73",x"81",x"c3"),
  1699 => (x"92",x"c2",x"9a",x"cf"),
  1700 => (x"30",x"72",x"48",x"c1"),
  1701 => (x"ba",x"ff",x"4a",x"70"),
  1702 => (x"98",x"69",x"48",x"72"),
  1703 => (x"87",x"db",x"79",x"70"),
  1704 => (x"b7",x"c4",x"49",x"73"),
  1705 => (x"ed",x"c1",x"91",x"29"),
  1706 => (x"4a",x"73",x"81",x"c3"),
  1707 => (x"92",x"c2",x"9a",x"cf"),
  1708 => (x"30",x"72",x"48",x"c3"),
  1709 => (x"69",x"48",x"4a",x"70"),
  1710 => (x"c1",x"79",x"70",x"b0"),
  1711 => (x"c0",x"48",x"e7",x"eb"),
  1712 => (x"e3",x"eb",x"c1",x"78"),
  1713 => (x"c2",x"78",x"c0",x"48"),
  1714 => (x"f9",x"49",x"c3",x"f8"),
  1715 => (x"4a",x"70",x"87",x"e3"),
  1716 => (x"03",x"aa",x"b7",x"c0"),
  1717 => (x"c0",x"87",x"dd",x"fd"),
  1718 => (x"26",x"87",x"c2",x"48"),
  1719 => (x"26",x"4c",x"26",x"4d"),
  1720 => (x"00",x"4f",x"26",x"4b"),
  1721 => (x"00",x"00",x"00",x"00"),
  1722 => (x"1e",x"00",x"00",x"00"),
  1723 => (x"fc",x"49",x"4a",x"71"),
  1724 => (x"4f",x"26",x"87",x"eb"),
  1725 => (x"72",x"4a",x"c0",x"1e"),
  1726 => (x"c1",x"91",x"c4",x"49"),
  1727 => (x"c0",x"81",x"c3",x"ed"),
  1728 => (x"d0",x"82",x"c1",x"79"),
  1729 => (x"ee",x"04",x"aa",x"b7"),
  1730 => (x"0e",x"4f",x"26",x"87"),
  1731 => (x"5d",x"5c",x"5b",x"5e"),
  1732 => (x"f8",x"4d",x"71",x"0e"),
  1733 => (x"4a",x"75",x"87",x"cb"),
  1734 => (x"92",x"2a",x"b7",x"c4"),
  1735 => (x"82",x"c3",x"ed",x"c1"),
  1736 => (x"9c",x"cf",x"4c",x"75"),
  1737 => (x"49",x"6a",x"94",x"c2"),
  1738 => (x"c3",x"2b",x"74",x"4b"),
  1739 => (x"74",x"48",x"c2",x"9b"),
  1740 => (x"ff",x"4c",x"70",x"30"),
  1741 => (x"71",x"48",x"74",x"bc"),
  1742 => (x"f7",x"7a",x"70",x"98"),
  1743 => (x"48",x"73",x"87",x"db"),
  1744 => (x"00",x"87",x"d8",x"fe"),
  1745 => (x"00",x"00",x"00",x"00"),
  1746 => (x"00",x"00",x"00",x"00"),
  1747 => (x"00",x"00",x"00",x"00"),
  1748 => (x"00",x"00",x"00",x"00"),
  1749 => (x"00",x"00",x"00",x"00"),
  1750 => (x"00",x"00",x"00",x"00"),
  1751 => (x"00",x"00",x"00",x"00"),
  1752 => (x"00",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"00",x"00",x"00",x"00"),
  1756 => (x"00",x"00",x"00",x"00"),
  1757 => (x"00",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"00",x"00"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"1e",x"00",x"00",x"00"),
  1761 => (x"c8",x"48",x"d0",x"ff"),
  1762 => (x"48",x"71",x"78",x"e1"),
  1763 => (x"78",x"08",x"d4",x"ff"),
  1764 => (x"ff",x"48",x"66",x"c4"),
  1765 => (x"26",x"78",x"08",x"d4"),
  1766 => (x"4a",x"71",x"1e",x"4f"),
  1767 => (x"1e",x"49",x"66",x"c4"),
  1768 => (x"de",x"ff",x"49",x"72"),
  1769 => (x"48",x"d0",x"ff",x"87"),
  1770 => (x"26",x"78",x"e0",x"c0"),
  1771 => (x"73",x"1e",x"4f",x"26"),
  1772 => (x"c8",x"4b",x"71",x"1e"),
  1773 => (x"73",x"1e",x"49",x"66"),
  1774 => (x"a2",x"e0",x"c1",x"4a"),
  1775 => (x"87",x"d9",x"ff",x"49"),
  1776 => (x"26",x"87",x"c4",x"26"),
  1777 => (x"26",x"4c",x"26",x"4d"),
  1778 => (x"1e",x"4f",x"26",x"4b"),
  1779 => (x"c3",x"4a",x"d4",x"ff"),
  1780 => (x"d0",x"ff",x"7a",x"ff"),
  1781 => (x"78",x"e1",x"c8",x"48"),
  1782 => (x"f8",x"c2",x"7a",x"de"),
  1783 => (x"49",x"7a",x"bf",x"cd"),
  1784 => (x"70",x"28",x"c8",x"48"),
  1785 => (x"d0",x"48",x"71",x"7a"),
  1786 => (x"71",x"7a",x"70",x"28"),
  1787 => (x"70",x"28",x"d8",x"48"),
  1788 => (x"48",x"d0",x"ff",x"7a"),
  1789 => (x"26",x"78",x"e0",x"c0"),
  1790 => (x"5b",x"5e",x"0e",x"4f"),
  1791 => (x"71",x"0e",x"5d",x"5c"),
  1792 => (x"cd",x"f8",x"c2",x"4c"),
  1793 => (x"74",x"4b",x"4d",x"bf"),
  1794 => (x"9b",x"66",x"d0",x"2b"),
  1795 => (x"66",x"d4",x"83",x"c1"),
  1796 => (x"87",x"c2",x"04",x"ab"),
  1797 => (x"4a",x"74",x"4b",x"c0"),
  1798 => (x"72",x"49",x"66",x"d0"),
  1799 => (x"75",x"b9",x"ff",x"31"),
  1800 => (x"72",x"48",x"73",x"99"),
  1801 => (x"48",x"4a",x"70",x"30"),
  1802 => (x"f8",x"c2",x"b0",x"71"),
  1803 => (x"da",x"fe",x"58",x"d1"),
  1804 => (x"26",x"4d",x"26",x"87"),
  1805 => (x"26",x"4b",x"26",x"4c"),
  1806 => (x"5b",x"5e",x"0e",x"4f"),
  1807 => (x"1e",x"0e",x"5d",x"5c"),
  1808 => (x"f8",x"c2",x"4c",x"71"),
  1809 => (x"4a",x"c0",x"4b",x"d1"),
  1810 => (x"fe",x"49",x"f4",x"c0"),
  1811 => (x"74",x"87",x"f6",x"d1"),
  1812 => (x"d1",x"f8",x"c2",x"1e"),
  1813 => (x"d8",x"ee",x"fe",x"49"),
  1814 => (x"70",x"86",x"c4",x"87"),
  1815 => (x"ea",x"c0",x"02",x"98"),
  1816 => (x"a6",x"1e",x"c4",x"87"),
  1817 => (x"f8",x"c2",x"1e",x"4d"),
  1818 => (x"f4",x"fe",x"49",x"d1"),
  1819 => (x"86",x"c8",x"87",x"c6"),
  1820 => (x"d6",x"02",x"98",x"70"),
  1821 => (x"c1",x"4a",x"75",x"87"),
  1822 => (x"c4",x"49",x"c1",x"f3"),
  1823 => (x"e9",x"cf",x"fe",x"4b"),
  1824 => (x"02",x"98",x"70",x"87"),
  1825 => (x"48",x"c0",x"87",x"ca"),
  1826 => (x"c0",x"87",x"ed",x"c0"),
  1827 => (x"87",x"e8",x"c0",x"48"),
  1828 => (x"c1",x"87",x"f3",x"c0"),
  1829 => (x"98",x"70",x"87",x"c4"),
  1830 => (x"c0",x"87",x"c8",x"02"),
  1831 => (x"98",x"70",x"87",x"fc"),
  1832 => (x"c2",x"87",x"f8",x"05"),
  1833 => (x"02",x"bf",x"f1",x"f8"),
  1834 => (x"f8",x"c2",x"87",x"cc"),
  1835 => (x"f8",x"c2",x"48",x"cd"),
  1836 => (x"fc",x"78",x"bf",x"f1"),
  1837 => (x"48",x"c1",x"87",x"d5"),
  1838 => (x"26",x"4d",x"26",x"26"),
  1839 => (x"26",x"4b",x"26",x"4c"),
  1840 => (x"52",x"41",x"5b",x"4f"),
  1841 => (x"c0",x"1e",x"00",x"43"),
  1842 => (x"d1",x"f8",x"c2",x"1e"),
  1843 => (x"fc",x"f0",x"fe",x"49"),
  1844 => (x"e9",x"f8",x"c2",x"87"),
  1845 => (x"26",x"78",x"c0",x"48"),
  1846 => (x"5e",x"0e",x"4f",x"26"),
  1847 => (x"0e",x"5d",x"5c",x"5b"),
  1848 => (x"a6",x"c4",x"86",x"f4"),
  1849 => (x"c2",x"78",x"c0",x"48"),
  1850 => (x"48",x"bf",x"e9",x"f8"),
  1851 => (x"03",x"a8",x"b7",x"c3"),
  1852 => (x"f8",x"c2",x"87",x"d1"),
  1853 => (x"c1",x"48",x"bf",x"e9"),
  1854 => (x"ed",x"f8",x"c2",x"80"),
  1855 => (x"48",x"fb",x"c0",x"58"),
  1856 => (x"c2",x"87",x"e2",x"c6"),
  1857 => (x"fe",x"49",x"d1",x"f8"),
  1858 => (x"70",x"87",x"fd",x"f5"),
  1859 => (x"e9",x"f8",x"c2",x"4c"),
  1860 => (x"8a",x"c3",x"4a",x"bf"),
  1861 => (x"c1",x"87",x"d8",x"02"),
  1862 => (x"cb",x"c5",x"02",x"8a"),
  1863 => (x"c2",x"02",x"8a",x"87"),
  1864 => (x"02",x"8a",x"87",x"f6"),
  1865 => (x"8a",x"87",x"cd",x"c1"),
  1866 => (x"87",x"e2",x"c3",x"02"),
  1867 => (x"c0",x"87",x"e1",x"c5"),
  1868 => (x"c4",x"4a",x"75",x"4d"),
  1869 => (x"c3",x"fb",x"c1",x"92"),
  1870 => (x"e5",x"f8",x"c2",x"82"),
  1871 => (x"70",x"80",x"75",x"48"),
  1872 => (x"bf",x"97",x"6e",x"7e"),
  1873 => (x"6e",x"4b",x"49",x"4b"),
  1874 => (x"50",x"a3",x"c1",x"48"),
  1875 => (x"48",x"11",x"81",x"6a"),
  1876 => (x"70",x"58",x"a6",x"cc"),
  1877 => (x"87",x"c4",x"02",x"ac"),
  1878 => (x"50",x"c0",x"48",x"6e"),
  1879 => (x"c7",x"05",x"66",x"c8"),
  1880 => (x"e9",x"f8",x"c2",x"87"),
  1881 => (x"78",x"a5",x"c4",x"48"),
  1882 => (x"b7",x"c4",x"85",x"c1"),
  1883 => (x"c0",x"ff",x"04",x"ad"),
  1884 => (x"87",x"dc",x"c4",x"87"),
  1885 => (x"bf",x"f5",x"f8",x"c2"),
  1886 => (x"a8",x"b7",x"c8",x"48"),
  1887 => (x"ca",x"87",x"d1",x"01"),
  1888 => (x"87",x"cc",x"02",x"ac"),
  1889 => (x"c7",x"02",x"ac",x"cd"),
  1890 => (x"ac",x"b7",x"c0",x"87"),
  1891 => (x"87",x"f3",x"c0",x"03"),
  1892 => (x"bf",x"f5",x"f8",x"c2"),
  1893 => (x"ab",x"b7",x"c8",x"4b"),
  1894 => (x"c2",x"87",x"d2",x"03"),
  1895 => (x"73",x"49",x"f9",x"f8"),
  1896 => (x"51",x"e0",x"c0",x"81"),
  1897 => (x"b7",x"c8",x"83",x"c1"),
  1898 => (x"ee",x"ff",x"04",x"ab"),
  1899 => (x"c1",x"f9",x"c2",x"87"),
  1900 => (x"50",x"d2",x"c1",x"48"),
  1901 => (x"c1",x"50",x"cf",x"c1"),
  1902 => (x"50",x"c0",x"50",x"cd"),
  1903 => (x"78",x"c3",x"80",x"e4"),
  1904 => (x"c2",x"87",x"cd",x"c3"),
  1905 => (x"49",x"bf",x"f5",x"f8"),
  1906 => (x"c2",x"80",x"c1",x"48"),
  1907 => (x"48",x"58",x"f9",x"f8"),
  1908 => (x"74",x"81",x"a0",x"c4"),
  1909 => (x"87",x"f8",x"c2",x"51"),
  1910 => (x"ac",x"b7",x"f0",x"c0"),
  1911 => (x"c0",x"87",x"da",x"04"),
  1912 => (x"01",x"ac",x"b7",x"f9"),
  1913 => (x"f8",x"c2",x"87",x"d3"),
  1914 => (x"ca",x"49",x"bf",x"ed"),
  1915 => (x"c0",x"4a",x"74",x"91"),
  1916 => (x"f8",x"c2",x"8a",x"f0"),
  1917 => (x"a1",x"72",x"48",x"ed"),
  1918 => (x"02",x"ac",x"ca",x"78"),
  1919 => (x"cd",x"87",x"c6",x"c0"),
  1920 => (x"cb",x"c2",x"05",x"ac"),
  1921 => (x"e9",x"f8",x"c2",x"87"),
  1922 => (x"c2",x"78",x"c3",x"48"),
  1923 => (x"f0",x"c0",x"87",x"c2"),
  1924 => (x"db",x"04",x"ac",x"b7"),
  1925 => (x"b7",x"f9",x"c0",x"87"),
  1926 => (x"d3",x"c0",x"01",x"ac"),
  1927 => (x"f1",x"f8",x"c2",x"87"),
  1928 => (x"91",x"d0",x"49",x"bf"),
  1929 => (x"f0",x"c0",x"4a",x"74"),
  1930 => (x"f1",x"f8",x"c2",x"8a"),
  1931 => (x"78",x"a1",x"72",x"48"),
  1932 => (x"ac",x"b7",x"c1",x"c1"),
  1933 => (x"87",x"db",x"c0",x"04"),
  1934 => (x"ac",x"b7",x"c6",x"c1"),
  1935 => (x"87",x"d3",x"c0",x"01"),
  1936 => (x"bf",x"f1",x"f8",x"c2"),
  1937 => (x"74",x"91",x"d0",x"49"),
  1938 => (x"8a",x"f7",x"c0",x"4a"),
  1939 => (x"48",x"f1",x"f8",x"c2"),
  1940 => (x"ca",x"78",x"a1",x"72"),
  1941 => (x"c6",x"c0",x"02",x"ac"),
  1942 => (x"05",x"ac",x"cd",x"87"),
  1943 => (x"c2",x"87",x"f1",x"c0"),
  1944 => (x"c3",x"48",x"e9",x"f8"),
  1945 => (x"87",x"e8",x"c0",x"78"),
  1946 => (x"05",x"ac",x"e2",x"c0"),
  1947 => (x"c4",x"87",x"c9",x"c0"),
  1948 => (x"fb",x"c0",x"48",x"a6"),
  1949 => (x"87",x"d8",x"c0",x"78"),
  1950 => (x"c0",x"02",x"ac",x"ca"),
  1951 => (x"ac",x"cd",x"87",x"c6"),
  1952 => (x"87",x"c9",x"c0",x"05"),
  1953 => (x"48",x"e9",x"f8",x"c2"),
  1954 => (x"c3",x"c0",x"78",x"c3"),
  1955 => (x"5c",x"a6",x"c8",x"87"),
  1956 => (x"03",x"ac",x"b7",x"c0"),
  1957 => (x"48",x"87",x"c4",x"c0"),
  1958 => (x"c4",x"87",x"ca",x"c0"),
  1959 => (x"c6",x"f9",x"02",x"66"),
  1960 => (x"ff",x"c3",x"48",x"87"),
  1961 => (x"f8",x"8e",x"f4",x"99"),
  1962 => (x"4f",x"43",x"87",x"cf"),
  1963 => (x"00",x"3d",x"46",x"4e"),
  1964 => (x"00",x"44",x"4f",x"4d"),
  1965 => (x"45",x"4d",x"41",x"4e"),
  1966 => (x"46",x"45",x"44",x"00"),
  1967 => (x"54",x"4c",x"55",x"41"),
  1968 => (x"aa",x"00",x"30",x"3d"),
  1969 => (x"b0",x"00",x"00",x"1e"),
  1970 => (x"b4",x"00",x"00",x"1e"),
  1971 => (x"b9",x"00",x"00",x"1e"),
  1972 => (x"1e",x"00",x"00",x"1e"),
  1973 => (x"c8",x"48",x"d0",x"ff"),
  1974 => (x"48",x"71",x"78",x"c9"),
  1975 => (x"78",x"08",x"d4",x"ff"),
  1976 => (x"71",x"1e",x"4f",x"26"),
  1977 => (x"87",x"eb",x"49",x"4a"),
  1978 => (x"c8",x"48",x"d0",x"ff"),
  1979 => (x"1e",x"4f",x"26",x"78"),
  1980 => (x"4b",x"71",x"1e",x"73"),
  1981 => (x"bf",x"d1",x"f9",x"c2"),
  1982 => (x"c2",x"87",x"c3",x"02"),
  1983 => (x"d0",x"ff",x"87",x"eb"),
  1984 => (x"78",x"c9",x"c8",x"48"),
  1985 => (x"e0",x"c0",x"49",x"73"),
  1986 => (x"48",x"d4",x"ff",x"b1"),
  1987 => (x"f9",x"c2",x"78",x"71"),
  1988 => (x"78",x"c0",x"48",x"c5"),
  1989 => (x"c5",x"02",x"66",x"c8"),
  1990 => (x"49",x"ff",x"c3",x"87"),
  1991 => (x"49",x"c0",x"87",x"c2"),
  1992 => (x"59",x"cd",x"f9",x"c2"),
  1993 => (x"c6",x"02",x"66",x"cc"),
  1994 => (x"d5",x"d5",x"c5",x"87"),
  1995 => (x"cf",x"87",x"c4",x"4a"),
  1996 => (x"c2",x"4a",x"ff",x"ff"),
  1997 => (x"c2",x"5a",x"d1",x"f9"),
  1998 => (x"c1",x"48",x"d1",x"f9"),
  1999 => (x"26",x"87",x"c4",x"78"),
  2000 => (x"26",x"4c",x"26",x"4d"),
  2001 => (x"0e",x"4f",x"26",x"4b"),
  2002 => (x"5d",x"5c",x"5b",x"5e"),
  2003 => (x"c2",x"4a",x"71",x"0e"),
  2004 => (x"4c",x"bf",x"cd",x"f9"),
  2005 => (x"cb",x"02",x"9a",x"72"),
  2006 => (x"91",x"c8",x"49",x"87"),
  2007 => (x"4b",x"e5",x"fb",x"c1"),
  2008 => (x"87",x"c4",x"83",x"71"),
  2009 => (x"4b",x"e5",x"ff",x"c1"),
  2010 => (x"49",x"13",x"4d",x"c0"),
  2011 => (x"f9",x"c2",x"99",x"74"),
  2012 => (x"ff",x"b9",x"bf",x"c9"),
  2013 => (x"78",x"71",x"48",x"d4"),
  2014 => (x"85",x"2c",x"b7",x"c1"),
  2015 => (x"04",x"ad",x"b7",x"c8"),
  2016 => (x"f9",x"c2",x"87",x"e8"),
  2017 => (x"c8",x"48",x"bf",x"c5"),
  2018 => (x"c9",x"f9",x"c2",x"80"),
  2019 => (x"87",x"ef",x"fe",x"58"),
  2020 => (x"71",x"1e",x"73",x"1e"),
  2021 => (x"9a",x"4a",x"13",x"4b"),
  2022 => (x"72",x"87",x"cb",x"02"),
  2023 => (x"87",x"e7",x"fe",x"49"),
  2024 => (x"05",x"9a",x"4a",x"13"),
  2025 => (x"da",x"fe",x"87",x"f5"),
  2026 => (x"f9",x"c2",x"1e",x"87"),
  2027 => (x"c2",x"49",x"bf",x"c5"),
  2028 => (x"c1",x"48",x"c5",x"f9"),
  2029 => (x"c0",x"c4",x"78",x"a1"),
  2030 => (x"db",x"03",x"a9",x"b7"),
  2031 => (x"48",x"d4",x"ff",x"87"),
  2032 => (x"bf",x"c9",x"f9",x"c2"),
  2033 => (x"c5",x"f9",x"c2",x"78"),
  2034 => (x"f9",x"c2",x"49",x"bf"),
  2035 => (x"a1",x"c1",x"48",x"c5"),
  2036 => (x"b7",x"c0",x"c4",x"78"),
  2037 => (x"87",x"e5",x"04",x"a9"),
  2038 => (x"c8",x"48",x"d0",x"ff"),
  2039 => (x"d1",x"f9",x"c2",x"78"),
  2040 => (x"26",x"78",x"c0",x"48"),
  2041 => (x"00",x"00",x"00",x"4f"),
  2042 => (x"00",x"00",x"00",x"00"),
  2043 => (x"00",x"00",x"00",x"00"),
  2044 => (x"00",x"00",x"5f",x"5f"),
  2045 => (x"03",x"03",x"00",x"00"),
  2046 => (x"00",x"03",x"03",x"00"),
  2047 => (x"7f",x"7f",x"14",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

