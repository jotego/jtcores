
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"14",x"7f",x"7f",x"14"),
     1 => (x"2e",x"24",x"00",x"00"),
     2 => (x"12",x"3a",x"6b",x"6b"),
     3 => (x"36",x"6a",x"4c",x"00"),
     4 => (x"32",x"56",x"6c",x"18"),
     5 => (x"4f",x"7e",x"30",x"00"),
     6 => (x"68",x"3a",x"77",x"59"),
     7 => (x"04",x"00",x"00",x"40"),
     8 => (x"00",x"00",x"03",x"07"),
     9 => (x"1c",x"00",x"00",x"00"),
    10 => (x"00",x"41",x"63",x"3e"),
    11 => (x"41",x"00",x"00",x"00"),
    12 => (x"00",x"1c",x"3e",x"63"),
    13 => (x"3e",x"2a",x"08",x"00"),
    14 => (x"2a",x"3e",x"1c",x"1c"),
    15 => (x"08",x"08",x"00",x"08"),
    16 => (x"08",x"08",x"3e",x"3e"),
    17 => (x"80",x"00",x"00",x"00"),
    18 => (x"00",x"00",x"60",x"e0"),
    19 => (x"08",x"08",x"00",x"00"),
    20 => (x"08",x"08",x"08",x"08"),
    21 => (x"00",x"00",x"00",x"00"),
    22 => (x"00",x"00",x"60",x"60"),
    23 => (x"30",x"60",x"40",x"00"),
    24 => (x"03",x"06",x"0c",x"18"),
    25 => (x"7f",x"3e",x"00",x"01"),
    26 => (x"3e",x"7f",x"4d",x"59"),
    27 => (x"06",x"04",x"00",x"00"),
    28 => (x"00",x"00",x"7f",x"7f"),
    29 => (x"63",x"42",x"00",x"00"),
    30 => (x"46",x"4f",x"59",x"71"),
    31 => (x"63",x"22",x"00",x"00"),
    32 => (x"36",x"7f",x"49",x"49"),
    33 => (x"16",x"1c",x"18",x"00"),
    34 => (x"10",x"7f",x"7f",x"13"),
    35 => (x"67",x"27",x"00",x"00"),
    36 => (x"39",x"7d",x"45",x"45"),
    37 => (x"7e",x"3c",x"00",x"00"),
    38 => (x"30",x"79",x"49",x"4b"),
    39 => (x"01",x"01",x"00",x"00"),
    40 => (x"07",x"0f",x"79",x"71"),
    41 => (x"7f",x"36",x"00",x"00"),
    42 => (x"36",x"7f",x"49",x"49"),
    43 => (x"4f",x"06",x"00",x"00"),
    44 => (x"1e",x"3f",x"69",x"49"),
    45 => (x"00",x"00",x"00",x"00"),
    46 => (x"00",x"00",x"66",x"66"),
    47 => (x"80",x"00",x"00",x"00"),
    48 => (x"00",x"00",x"66",x"e6"),
    49 => (x"08",x"08",x"00",x"00"),
    50 => (x"22",x"22",x"14",x"14"),
    51 => (x"14",x"14",x"00",x"00"),
    52 => (x"14",x"14",x"14",x"14"),
    53 => (x"22",x"22",x"00",x"00"),
    54 => (x"08",x"08",x"14",x"14"),
    55 => (x"03",x"02",x"00",x"00"),
    56 => (x"06",x"0f",x"59",x"51"),
    57 => (x"41",x"7f",x"3e",x"00"),
    58 => (x"1e",x"1f",x"55",x"5d"),
    59 => (x"7f",x"7e",x"00",x"00"),
    60 => (x"7e",x"7f",x"09",x"09"),
    61 => (x"7f",x"7f",x"00",x"00"),
    62 => (x"36",x"7f",x"49",x"49"),
    63 => (x"3e",x"1c",x"00",x"00"),
    64 => (x"41",x"41",x"41",x"63"),
    65 => (x"7f",x"7f",x"00",x"00"),
    66 => (x"1c",x"3e",x"63",x"41"),
    67 => (x"7f",x"7f",x"00",x"00"),
    68 => (x"41",x"41",x"49",x"49"),
    69 => (x"7f",x"7f",x"00",x"00"),
    70 => (x"01",x"01",x"09",x"09"),
    71 => (x"7f",x"3e",x"00",x"00"),
    72 => (x"7a",x"7b",x"49",x"41"),
    73 => (x"7f",x"7f",x"00",x"00"),
    74 => (x"7f",x"7f",x"08",x"08"),
    75 => (x"41",x"00",x"00",x"00"),
    76 => (x"00",x"41",x"7f",x"7f"),
    77 => (x"60",x"20",x"00",x"00"),
    78 => (x"3f",x"7f",x"40",x"40"),
    79 => (x"08",x"7f",x"7f",x"00"),
    80 => (x"41",x"63",x"36",x"1c"),
    81 => (x"7f",x"7f",x"00",x"00"),
    82 => (x"40",x"40",x"40",x"40"),
    83 => (x"06",x"7f",x"7f",x"00"),
    84 => (x"7f",x"7f",x"06",x"0c"),
    85 => (x"06",x"7f",x"7f",x"00"),
    86 => (x"7f",x"7f",x"18",x"0c"),
    87 => (x"7f",x"3e",x"00",x"00"),
    88 => (x"3e",x"7f",x"41",x"41"),
    89 => (x"7f",x"7f",x"00",x"00"),
    90 => (x"06",x"0f",x"09",x"09"),
    91 => (x"41",x"7f",x"3e",x"00"),
    92 => (x"40",x"7e",x"7f",x"61"),
    93 => (x"7f",x"7f",x"00",x"00"),
    94 => (x"66",x"7f",x"19",x"09"),
    95 => (x"6f",x"26",x"00",x"00"),
    96 => (x"32",x"7b",x"59",x"4d"),
    97 => (x"01",x"01",x"00",x"00"),
    98 => (x"01",x"01",x"7f",x"7f"),
    99 => (x"7f",x"3f",x"00",x"00"),
   100 => (x"3f",x"7f",x"40",x"40"),
   101 => (x"3f",x"0f",x"00",x"00"),
   102 => (x"0f",x"3f",x"70",x"70"),
   103 => (x"30",x"7f",x"7f",x"00"),
   104 => (x"7f",x"7f",x"30",x"18"),
   105 => (x"36",x"63",x"41",x"00"),
   106 => (x"63",x"36",x"1c",x"1c"),
   107 => (x"06",x"03",x"01",x"41"),
   108 => (x"03",x"06",x"7c",x"7c"),
   109 => (x"59",x"71",x"61",x"01"),
   110 => (x"41",x"43",x"47",x"4d"),
   111 => (x"7f",x"00",x"00",x"00"),
   112 => (x"00",x"41",x"41",x"7f"),
   113 => (x"06",x"03",x"01",x"00"),
   114 => (x"60",x"30",x"18",x"0c"),
   115 => (x"41",x"00",x"00",x"40"),
   116 => (x"00",x"7f",x"7f",x"41"),
   117 => (x"06",x"0c",x"08",x"00"),
   118 => (x"08",x"0c",x"06",x"03"),
   119 => (x"80",x"80",x"80",x"00"),
   120 => (x"80",x"80",x"80",x"80"),
   121 => (x"00",x"00",x"00",x"00"),
   122 => (x"00",x"04",x"07",x"03"),
   123 => (x"74",x"20",x"00",x"00"),
   124 => (x"78",x"7c",x"54",x"54"),
   125 => (x"7f",x"7f",x"00",x"00"),
   126 => (x"38",x"7c",x"44",x"44"),
   127 => (x"7c",x"38",x"00",x"00"),
   128 => (x"00",x"44",x"44",x"44"),
   129 => (x"7c",x"38",x"00",x"00"),
   130 => (x"7f",x"7f",x"44",x"44"),
   131 => (x"7c",x"38",x"00",x"00"),
   132 => (x"18",x"5c",x"54",x"54"),
   133 => (x"7e",x"04",x"00",x"00"),
   134 => (x"00",x"05",x"05",x"7f"),
   135 => (x"bc",x"18",x"00",x"00"),
   136 => (x"7c",x"fc",x"a4",x"a4"),
   137 => (x"7f",x"7f",x"00",x"00"),
   138 => (x"78",x"7c",x"04",x"04"),
   139 => (x"00",x"00",x"00",x"00"),
   140 => (x"00",x"40",x"7d",x"3d"),
   141 => (x"80",x"80",x"00",x"00"),
   142 => (x"00",x"7d",x"fd",x"80"),
   143 => (x"7f",x"7f",x"00",x"00"),
   144 => (x"44",x"6c",x"38",x"10"),
   145 => (x"00",x"00",x"00",x"00"),
   146 => (x"00",x"40",x"7f",x"3f"),
   147 => (x"0c",x"7c",x"7c",x"00"),
   148 => (x"78",x"7c",x"0c",x"18"),
   149 => (x"7c",x"7c",x"00",x"00"),
   150 => (x"78",x"7c",x"04",x"04"),
   151 => (x"7c",x"38",x"00",x"00"),
   152 => (x"38",x"7c",x"44",x"44"),
   153 => (x"fc",x"fc",x"00",x"00"),
   154 => (x"18",x"3c",x"24",x"24"),
   155 => (x"3c",x"18",x"00",x"00"),
   156 => (x"fc",x"fc",x"24",x"24"),
   157 => (x"7c",x"7c",x"00",x"00"),
   158 => (x"08",x"0c",x"04",x"04"),
   159 => (x"5c",x"48",x"00",x"00"),
   160 => (x"20",x"74",x"54",x"54"),
   161 => (x"3f",x"04",x"00",x"00"),
   162 => (x"00",x"44",x"44",x"7f"),
   163 => (x"7c",x"3c",x"00",x"00"),
   164 => (x"7c",x"7c",x"40",x"40"),
   165 => (x"3c",x"1c",x"00",x"00"),
   166 => (x"1c",x"3c",x"60",x"60"),
   167 => (x"60",x"7c",x"3c",x"00"),
   168 => (x"3c",x"7c",x"60",x"30"),
   169 => (x"38",x"6c",x"44",x"00"),
   170 => (x"44",x"6c",x"38",x"10"),
   171 => (x"bc",x"1c",x"00",x"00"),
   172 => (x"1c",x"3c",x"60",x"e0"),
   173 => (x"64",x"44",x"00",x"00"),
   174 => (x"44",x"4c",x"5c",x"74"),
   175 => (x"08",x"08",x"00",x"00"),
   176 => (x"41",x"41",x"77",x"3e"),
   177 => (x"00",x"00",x"00",x"00"),
   178 => (x"00",x"00",x"7f",x"7f"),
   179 => (x"41",x"41",x"00",x"00"),
   180 => (x"08",x"08",x"3e",x"77"),
   181 => (x"01",x"01",x"02",x"00"),
   182 => (x"01",x"02",x"02",x"03"),
   183 => (x"7f",x"7f",x"7f",x"00"),
   184 => (x"7f",x"7f",x"7f",x"7f"),
   185 => (x"1c",x"08",x"08",x"00"),
   186 => (x"7f",x"3e",x"3e",x"1c"),
   187 => (x"3e",x"7f",x"7f",x"7f"),
   188 => (x"08",x"1c",x"1c",x"3e"),
   189 => (x"18",x"10",x"00",x"08"),
   190 => (x"10",x"18",x"7c",x"7c"),
   191 => (x"30",x"10",x"00",x"00"),
   192 => (x"10",x"30",x"7c",x"7c"),
   193 => (x"60",x"30",x"10",x"00"),
   194 => (x"06",x"1e",x"78",x"60"),
   195 => (x"3c",x"66",x"42",x"00"),
   196 => (x"42",x"66",x"3c",x"18"),
   197 => (x"6a",x"38",x"78",x"00"),
   198 => (x"38",x"6c",x"c6",x"c2"),
   199 => (x"00",x"00",x"60",x"00"),
   200 => (x"60",x"00",x"00",x"60"),
   201 => (x"5b",x"5e",x"0e",x"00"),
   202 => (x"1e",x"0e",x"5d",x"5c"),
   203 => (x"f9",x"c2",x"4c",x"71"),
   204 => (x"c0",x"4d",x"bf",x"e2"),
   205 => (x"74",x"1e",x"c0",x"4b"),
   206 => (x"87",x"c7",x"02",x"ab"),
   207 => (x"c0",x"48",x"a6",x"c4"),
   208 => (x"c4",x"87",x"c5",x"78"),
   209 => (x"78",x"c1",x"48",x"a6"),
   210 => (x"73",x"1e",x"66",x"c4"),
   211 => (x"87",x"df",x"ee",x"49"),
   212 => (x"e0",x"c0",x"86",x"c8"),
   213 => (x"87",x"ef",x"ef",x"49"),
   214 => (x"6a",x"4a",x"a5",x"c4"),
   215 => (x"87",x"f0",x"f0",x"49"),
   216 => (x"cb",x"87",x"c6",x"f1"),
   217 => (x"c8",x"83",x"c1",x"85"),
   218 => (x"ff",x"04",x"ab",x"b7"),
   219 => (x"26",x"26",x"87",x"c7"),
   220 => (x"26",x"4c",x"26",x"4d"),
   221 => (x"1e",x"4f",x"26",x"4b"),
   222 => (x"f9",x"c2",x"4a",x"71"),
   223 => (x"f9",x"c2",x"5a",x"e6"),
   224 => (x"78",x"c7",x"48",x"e6"),
   225 => (x"87",x"dd",x"fe",x"49"),
   226 => (x"73",x"1e",x"4f",x"26"),
   227 => (x"c0",x"4a",x"71",x"1e"),
   228 => (x"d3",x"03",x"aa",x"b7"),
   229 => (x"ea",x"db",x"c2",x"87"),
   230 => (x"87",x"c4",x"05",x"bf"),
   231 => (x"87",x"c2",x"4b",x"c1"),
   232 => (x"db",x"c2",x"4b",x"c0"),
   233 => (x"87",x"c4",x"5b",x"ee"),
   234 => (x"5a",x"ee",x"db",x"c2"),
   235 => (x"bf",x"ea",x"db",x"c2"),
   236 => (x"c1",x"9a",x"c1",x"4a"),
   237 => (x"ec",x"49",x"a2",x"c0"),
   238 => (x"48",x"fc",x"87",x"e8"),
   239 => (x"bf",x"ea",x"db",x"c2"),
   240 => (x"87",x"ef",x"fe",x"78"),
   241 => (x"c4",x"4a",x"71",x"1e"),
   242 => (x"49",x"72",x"1e",x"66"),
   243 => (x"87",x"de",x"df",x"ff"),
   244 => (x"1e",x"4f",x"26",x"26"),
   245 => (x"bf",x"ea",x"db",x"c2"),
   246 => (x"ce",x"dc",x"ff",x"49"),
   247 => (x"da",x"f9",x"c2",x"87"),
   248 => (x"78",x"bf",x"e8",x"48"),
   249 => (x"48",x"d6",x"f9",x"c2"),
   250 => (x"c2",x"78",x"bf",x"ec"),
   251 => (x"4a",x"bf",x"da",x"f9"),
   252 => (x"99",x"ff",x"c3",x"49"),
   253 => (x"72",x"2a",x"b7",x"c8"),
   254 => (x"c2",x"b0",x"71",x"48"),
   255 => (x"26",x"58",x"e2",x"f9"),
   256 => (x"5b",x"5e",x"0e",x"4f"),
   257 => (x"71",x"0e",x"5d",x"5c"),
   258 => (x"87",x"c7",x"ff",x"4b"),
   259 => (x"48",x"d5",x"f9",x"c2"),
   260 => (x"49",x"73",x"50",x"c0"),
   261 => (x"87",x"f3",x"db",x"ff"),
   262 => (x"c2",x"4c",x"49",x"70"),
   263 => (x"49",x"ee",x"cb",x"9c"),
   264 => (x"70",x"87",x"cf",x"cb"),
   265 => (x"f9",x"c2",x"4d",x"49"),
   266 => (x"05",x"bf",x"97",x"d5"),
   267 => (x"d0",x"87",x"e4",x"c1"),
   268 => (x"f9",x"c2",x"49",x"66"),
   269 => (x"05",x"99",x"bf",x"de"),
   270 => (x"66",x"d4",x"87",x"d7"),
   271 => (x"d6",x"f9",x"c2",x"49"),
   272 => (x"cc",x"05",x"99",x"bf"),
   273 => (x"ff",x"49",x"73",x"87"),
   274 => (x"70",x"87",x"c0",x"db"),
   275 => (x"c2",x"c1",x"02",x"98"),
   276 => (x"fd",x"4c",x"c1",x"87"),
   277 => (x"49",x"75",x"87",x"fd"),
   278 => (x"70",x"87",x"e3",x"ca"),
   279 => (x"87",x"c6",x"02",x"98"),
   280 => (x"48",x"d5",x"f9",x"c2"),
   281 => (x"f9",x"c2",x"50",x"c1"),
   282 => (x"05",x"bf",x"97",x"d5"),
   283 => (x"c2",x"87",x"e4",x"c0"),
   284 => (x"49",x"bf",x"de",x"f9"),
   285 => (x"05",x"99",x"66",x"d0"),
   286 => (x"c2",x"87",x"d6",x"ff"),
   287 => (x"49",x"bf",x"d6",x"f9"),
   288 => (x"05",x"99",x"66",x"d4"),
   289 => (x"73",x"87",x"ca",x"ff"),
   290 => (x"fe",x"d9",x"ff",x"49"),
   291 => (x"05",x"98",x"70",x"87"),
   292 => (x"74",x"87",x"fe",x"fe"),
   293 => (x"87",x"d7",x"fb",x"48"),
   294 => (x"5c",x"5b",x"5e",x"0e"),
   295 => (x"86",x"f4",x"0e",x"5d"),
   296 => (x"ec",x"4c",x"4d",x"c0"),
   297 => (x"a6",x"c4",x"7e",x"bf"),
   298 => (x"e2",x"f9",x"c2",x"48"),
   299 => (x"1e",x"c1",x"78",x"bf"),
   300 => (x"49",x"c7",x"1e",x"c0"),
   301 => (x"c8",x"87",x"ca",x"fd"),
   302 => (x"02",x"98",x"70",x"86"),
   303 => (x"49",x"ff",x"87",x"ce"),
   304 => (x"c1",x"87",x"c7",x"fb"),
   305 => (x"d9",x"ff",x"49",x"da"),
   306 => (x"4d",x"c1",x"87",x"c1"),
   307 => (x"97",x"d5",x"f9",x"c2"),
   308 => (x"87",x"c3",x"02",x"bf"),
   309 => (x"c2",x"87",x"f9",x"cd"),
   310 => (x"4b",x"bf",x"da",x"f9"),
   311 => (x"bf",x"ea",x"db",x"c2"),
   312 => (x"87",x"eb",x"c0",x"05"),
   313 => (x"ff",x"49",x"fd",x"c3"),
   314 => (x"c3",x"87",x"e0",x"d8"),
   315 => (x"d8",x"ff",x"49",x"fa"),
   316 => (x"49",x"73",x"87",x"d9"),
   317 => (x"71",x"99",x"ff",x"c3"),
   318 => (x"fb",x"49",x"c0",x"1e"),
   319 => (x"49",x"73",x"87",x"c6"),
   320 => (x"71",x"29",x"b7",x"c8"),
   321 => (x"fa",x"49",x"c1",x"1e"),
   322 => (x"86",x"c8",x"87",x"fa"),
   323 => (x"c2",x"87",x"c1",x"c6"),
   324 => (x"4b",x"bf",x"de",x"f9"),
   325 => (x"87",x"dd",x"02",x"9b"),
   326 => (x"bf",x"e6",x"db",x"c2"),
   327 => (x"87",x"de",x"c7",x"49"),
   328 => (x"c4",x"05",x"98",x"70"),
   329 => (x"d2",x"4b",x"c0",x"87"),
   330 => (x"49",x"e0",x"c2",x"87"),
   331 => (x"c2",x"87",x"c3",x"c7"),
   332 => (x"c6",x"58",x"ea",x"db"),
   333 => (x"e6",x"db",x"c2",x"87"),
   334 => (x"73",x"78",x"c0",x"48"),
   335 => (x"05",x"99",x"c2",x"49"),
   336 => (x"eb",x"c3",x"87",x"ce"),
   337 => (x"c2",x"d7",x"ff",x"49"),
   338 => (x"c2",x"49",x"70",x"87"),
   339 => (x"87",x"c2",x"02",x"99"),
   340 => (x"49",x"73",x"4c",x"fb"),
   341 => (x"ce",x"05",x"99",x"c1"),
   342 => (x"49",x"f4",x"c3",x"87"),
   343 => (x"87",x"eb",x"d6",x"ff"),
   344 => (x"99",x"c2",x"49",x"70"),
   345 => (x"fa",x"87",x"c2",x"02"),
   346 => (x"c8",x"49",x"73",x"4c"),
   347 => (x"87",x"ce",x"05",x"99"),
   348 => (x"ff",x"49",x"f5",x"c3"),
   349 => (x"70",x"87",x"d4",x"d6"),
   350 => (x"02",x"99",x"c2",x"49"),
   351 => (x"f9",x"c2",x"87",x"d5"),
   352 => (x"ca",x"02",x"bf",x"e6"),
   353 => (x"88",x"c1",x"48",x"87"),
   354 => (x"58",x"ea",x"f9",x"c2"),
   355 => (x"ff",x"87",x"c2",x"c0"),
   356 => (x"73",x"4d",x"c1",x"4c"),
   357 => (x"05",x"99",x"c4",x"49"),
   358 => (x"f2",x"c3",x"87",x"ce"),
   359 => (x"ea",x"d5",x"ff",x"49"),
   360 => (x"c2",x"49",x"70",x"87"),
   361 => (x"87",x"dc",x"02",x"99"),
   362 => (x"bf",x"e6",x"f9",x"c2"),
   363 => (x"b7",x"c7",x"48",x"7e"),
   364 => (x"cb",x"c0",x"03",x"a8"),
   365 => (x"c1",x"48",x"6e",x"87"),
   366 => (x"ea",x"f9",x"c2",x"80"),
   367 => (x"87",x"c2",x"c0",x"58"),
   368 => (x"4d",x"c1",x"4c",x"fe"),
   369 => (x"ff",x"49",x"fd",x"c3"),
   370 => (x"70",x"87",x"c0",x"d5"),
   371 => (x"02",x"99",x"c2",x"49"),
   372 => (x"c2",x"87",x"d5",x"c0"),
   373 => (x"02",x"bf",x"e6",x"f9"),
   374 => (x"c2",x"87",x"c9",x"c0"),
   375 => (x"c0",x"48",x"e6",x"f9"),
   376 => (x"87",x"c2",x"c0",x"78"),
   377 => (x"4d",x"c1",x"4c",x"fd"),
   378 => (x"ff",x"49",x"fa",x"c3"),
   379 => (x"70",x"87",x"dc",x"d4"),
   380 => (x"02",x"99",x"c2",x"49"),
   381 => (x"c2",x"87",x"d9",x"c0"),
   382 => (x"48",x"bf",x"e6",x"f9"),
   383 => (x"03",x"a8",x"b7",x"c7"),
   384 => (x"c2",x"87",x"c9",x"c0"),
   385 => (x"c7",x"48",x"e6",x"f9"),
   386 => (x"87",x"c2",x"c0",x"78"),
   387 => (x"4d",x"c1",x"4c",x"fc"),
   388 => (x"03",x"ac",x"b7",x"c0"),
   389 => (x"c4",x"87",x"d1",x"c0"),
   390 => (x"d8",x"c1",x"4a",x"66"),
   391 => (x"c0",x"02",x"6a",x"82"),
   392 => (x"4b",x"6a",x"87",x"c6"),
   393 => (x"0f",x"73",x"49",x"74"),
   394 => (x"f0",x"c3",x"1e",x"c0"),
   395 => (x"49",x"da",x"c1",x"1e"),
   396 => (x"c8",x"87",x"ce",x"f7"),
   397 => (x"02",x"98",x"70",x"86"),
   398 => (x"c8",x"87",x"e2",x"c0"),
   399 => (x"f9",x"c2",x"48",x"a6"),
   400 => (x"c8",x"78",x"bf",x"e6"),
   401 => (x"91",x"cb",x"49",x"66"),
   402 => (x"71",x"48",x"66",x"c4"),
   403 => (x"6e",x"7e",x"70",x"80"),
   404 => (x"c8",x"c0",x"02",x"bf"),
   405 => (x"4b",x"bf",x"6e",x"87"),
   406 => (x"73",x"49",x"66",x"c8"),
   407 => (x"02",x"9d",x"75",x"0f"),
   408 => (x"c2",x"87",x"c8",x"c0"),
   409 => (x"49",x"bf",x"e6",x"f9"),
   410 => (x"c2",x"87",x"fa",x"f2"),
   411 => (x"02",x"bf",x"ee",x"db"),
   412 => (x"49",x"87",x"dd",x"c0"),
   413 => (x"70",x"87",x"c7",x"c2"),
   414 => (x"d3",x"c0",x"02",x"98"),
   415 => (x"e6",x"f9",x"c2",x"87"),
   416 => (x"e0",x"f2",x"49",x"bf"),
   417 => (x"f4",x"49",x"c0",x"87"),
   418 => (x"db",x"c2",x"87",x"c0"),
   419 => (x"78",x"c0",x"48",x"ee"),
   420 => (x"da",x"f3",x"8e",x"f4"),
   421 => (x"5b",x"5e",x"0e",x"87"),
   422 => (x"1e",x"0e",x"5d",x"5c"),
   423 => (x"f9",x"c2",x"4c",x"71"),
   424 => (x"c1",x"49",x"bf",x"e2"),
   425 => (x"c1",x"4d",x"a1",x"cd"),
   426 => (x"7e",x"69",x"81",x"d1"),
   427 => (x"cf",x"02",x"9c",x"74"),
   428 => (x"4b",x"a5",x"c4",x"87"),
   429 => (x"f9",x"c2",x"7b",x"74"),
   430 => (x"f2",x"49",x"bf",x"e2"),
   431 => (x"7b",x"6e",x"87",x"f9"),
   432 => (x"c4",x"05",x"9c",x"74"),
   433 => (x"c2",x"4b",x"c0",x"87"),
   434 => (x"73",x"4b",x"c1",x"87"),
   435 => (x"87",x"fa",x"f2",x"49"),
   436 => (x"c7",x"02",x"66",x"d4"),
   437 => (x"87",x"da",x"49",x"87"),
   438 => (x"87",x"c2",x"4a",x"70"),
   439 => (x"db",x"c2",x"4a",x"c0"),
   440 => (x"f2",x"26",x"5a",x"f2"),
   441 => (x"00",x"00",x"87",x"c9"),
   442 => (x"00",x"00",x"00",x"00"),
   443 => (x"00",x"00",x"00",x"00"),
   444 => (x"71",x"1e",x"00",x"00"),
   445 => (x"bf",x"c8",x"ff",x"4a"),
   446 => (x"48",x"a1",x"72",x"49"),
   447 => (x"ff",x"1e",x"4f",x"26"),
   448 => (x"fe",x"89",x"bf",x"c8"),
   449 => (x"c0",x"c0",x"c0",x"c0"),
   450 => (x"c4",x"01",x"a9",x"c0"),
   451 => (x"c2",x"4a",x"c0",x"87"),
   452 => (x"72",x"4a",x"c1",x"87"),
   453 => (x"0e",x"4f",x"26",x"48"),
   454 => (x"5d",x"5c",x"5b",x"5e"),
   455 => (x"4d",x"71",x"1e",x"0e"),
   456 => (x"75",x"4b",x"d4",x"ff"),
   457 => (x"ea",x"f9",x"c2",x"1e"),
   458 => (x"c4",x"c3",x"fe",x"49"),
   459 => (x"70",x"86",x"c4",x"87"),
   460 => (x"c3",x"02",x"6e",x"7e"),
   461 => (x"f9",x"c2",x"87",x"ff"),
   462 => (x"75",x"4c",x"bf",x"f2"),
   463 => (x"f4",x"dd",x"fe",x"49"),
   464 => (x"05",x"a8",x"de",x"87"),
   465 => (x"75",x"87",x"eb",x"c0"),
   466 => (x"ec",x"d3",x"ff",x"49"),
   467 => (x"02",x"98",x"70",x"87"),
   468 => (x"f8",x"c2",x"87",x"db"),
   469 => (x"c0",x"1e",x"bf",x"ed"),
   470 => (x"d0",x"ff",x"49",x"e1"),
   471 => (x"86",x"c4",x"87",x"fb"),
   472 => (x"48",x"cf",x"e1",x"c2"),
   473 => (x"f8",x"c2",x"50",x"c0"),
   474 => (x"ea",x"fe",x"49",x"f9"),
   475 => (x"c3",x"48",x"c1",x"87"),
   476 => (x"d0",x"ff",x"87",x"c5"),
   477 => (x"78",x"c5",x"c8",x"48"),
   478 => (x"c0",x"7b",x"d6",x"c1"),
   479 => (x"bf",x"97",x"6e",x"4a"),
   480 => (x"c1",x"48",x"6e",x"7b"),
   481 => (x"c1",x"7e",x"70",x"80"),
   482 => (x"b7",x"e0",x"c0",x"82"),
   483 => (x"ec",x"ff",x"04",x"aa"),
   484 => (x"48",x"d0",x"ff",x"87"),
   485 => (x"c5",x"c8",x"78",x"c4"),
   486 => (x"7b",x"d3",x"c1",x"78"),
   487 => (x"78",x"c4",x"7b",x"c1"),
   488 => (x"c1",x"02",x"9c",x"74"),
   489 => (x"e7",x"c2",x"87",x"fd"),
   490 => (x"c0",x"c8",x"7e",x"e6"),
   491 => (x"b7",x"c0",x"8c",x"4d"),
   492 => (x"87",x"c6",x"03",x"ac"),
   493 => (x"4d",x"a4",x"c0",x"c8"),
   494 => (x"f4",x"c2",x"4c",x"c0"),
   495 => (x"49",x"bf",x"97",x"d7"),
   496 => (x"d2",x"02",x"99",x"d0"),
   497 => (x"c2",x"1e",x"c0",x"87"),
   498 => (x"fe",x"49",x"ea",x"f9"),
   499 => (x"c4",x"87",x"f7",x"c3"),
   500 => (x"4a",x"49",x"70",x"86"),
   501 => (x"c2",x"87",x"ef",x"c0"),
   502 => (x"c2",x"1e",x"e6",x"e7"),
   503 => (x"fe",x"49",x"ea",x"f9"),
   504 => (x"c4",x"87",x"e3",x"c3"),
   505 => (x"4a",x"49",x"70",x"86"),
   506 => (x"c8",x"48",x"d0",x"ff"),
   507 => (x"d4",x"c1",x"78",x"c5"),
   508 => (x"bf",x"97",x"6e",x"7b"),
   509 => (x"c1",x"48",x"6e",x"7b"),
   510 => (x"c1",x"7e",x"70",x"80"),
   511 => (x"f0",x"ff",x"05",x"8d"),
   512 => (x"48",x"d0",x"ff",x"87"),
   513 => (x"9a",x"72",x"78",x"c4"),
   514 => (x"87",x"c5",x"c0",x"05"),
   515 => (x"e6",x"c0",x"48",x"c0"),
   516 => (x"c2",x"1e",x"c1",x"87"),
   517 => (x"fe",x"49",x"ea",x"f9"),
   518 => (x"c4",x"87",x"d1",x"c1"),
   519 => (x"05",x"9c",x"74",x"86"),
   520 => (x"ff",x"87",x"c3",x"fe"),
   521 => (x"c5",x"c8",x"48",x"d0"),
   522 => (x"7b",x"d3",x"c1",x"78"),
   523 => (x"78",x"c4",x"7b",x"c0"),
   524 => (x"c2",x"c0",x"48",x"c1"),
   525 => (x"26",x"48",x"c0",x"87"),
   526 => (x"4c",x"26",x"4d",x"26"),
   527 => (x"4f",x"26",x"4b",x"26"),
   528 => (x"c4",x"4a",x"71",x"1e"),
   529 => (x"87",x"c5",x"05",x"66"),
   530 => (x"ca",x"fb",x"49",x"72"),
   531 => (x"00",x"4f",x"26",x"87"),
   532 => (x"de",x"e2",x"c2",x"1e"),
   533 => (x"b9",x"c1",x"49",x"bf"),
   534 => (x"59",x"e2",x"e2",x"c2"),
   535 => (x"c3",x"48",x"d4",x"ff"),
   536 => (x"d0",x"ff",x"78",x"ff"),
   537 => (x"78",x"e1",x"c8",x"48"),
   538 => (x"c1",x"48",x"d4",x"ff"),
   539 => (x"71",x"31",x"c4",x"78"),
   540 => (x"48",x"d0",x"ff",x"78"),
   541 => (x"26",x"78",x"e0",x"c0"),
   542 => (x"e2",x"c2",x"1e",x"4f"),
   543 => (x"f9",x"c2",x"1e",x"d2"),
   544 => (x"fd",x"fd",x"49",x"ea"),
   545 => (x"86",x"c4",x"87",x"eb"),
   546 => (x"c3",x"02",x"98",x"70"),
   547 => (x"87",x"c0",x"ff",x"87"),
   548 => (x"35",x"31",x"4f",x"26"),
   549 => (x"20",x"5a",x"48",x"4b"),
   550 => (x"46",x"43",x"20",x"20"),
   551 => (x"00",x"00",x"00",x"47"),
   552 => (x"5e",x"0e",x"00",x"00"),
   553 => (x"0e",x"5d",x"5c",x"5b"),
   554 => (x"bf",x"d6",x"f9",x"c2"),
   555 => (x"cb",x"e4",x"c2",x"4a"),
   556 => (x"72",x"4c",x"49",x"bf"),
   557 => (x"ff",x"4d",x"71",x"bc"),
   558 => (x"c0",x"87",x"e6",x"c1"),
   559 => (x"d0",x"49",x"74",x"4b"),
   560 => (x"e7",x"c0",x"02",x"99"),
   561 => (x"48",x"d0",x"ff",x"87"),
   562 => (x"ff",x"78",x"e1",x"c8"),
   563 => (x"78",x"c5",x"48",x"d4"),
   564 => (x"99",x"d0",x"49",x"75"),
   565 => (x"c3",x"87",x"c3",x"02"),
   566 => (x"e6",x"c2",x"78",x"f0"),
   567 => (x"81",x"73",x"49",x"f7"),
   568 => (x"d4",x"ff",x"48",x"11"),
   569 => (x"d0",x"ff",x"78",x"08"),
   570 => (x"78",x"e0",x"c0",x"48"),
   571 => (x"83",x"2d",x"2c",x"c1"),
   572 => (x"ff",x"04",x"ab",x"c8"),
   573 => (x"c0",x"ff",x"87",x"c7"),
   574 => (x"e4",x"c2",x"87",x"df"),
   575 => (x"f9",x"c2",x"48",x"cb"),
   576 => (x"26",x"78",x"bf",x"d6"),
   577 => (x"26",x"4c",x"26",x"4d"),
   578 => (x"00",x"4f",x"26",x"4b"),
   579 => (x"1e",x"00",x"00",x"00"),
   580 => (x"4b",x"c0",x"1e",x"73"),
   581 => (x"48",x"cf",x"e1",x"c2"),
   582 => (x"1e",x"c8",x"50",x"de"),
   583 => (x"49",x"fe",x"f9",x"c2"),
   584 => (x"87",x"d0",x"d5",x"fe"),
   585 => (x"1e",x"72",x"86",x"c4"),
   586 => (x"48",x"c0",x"e6",x"c2"),
   587 => (x"49",x"c6",x"fa",x"c2"),
   588 => (x"20",x"4a",x"a1",x"c4"),
   589 => (x"05",x"aa",x"71",x"41"),
   590 => (x"4a",x"26",x"87",x"f9"),
   591 => (x"49",x"c4",x"e6",x"c2"),
   592 => (x"87",x"ce",x"f9",x"fd"),
   593 => (x"02",x"9a",x"4a",x"70"),
   594 => (x"fe",x"49",x"87",x"c5"),
   595 => (x"72",x"87",x"ef",x"c7"),
   596 => (x"d0",x"e6",x"c2",x"1e"),
   597 => (x"c6",x"fa",x"c2",x"48"),
   598 => (x"4a",x"a1",x"c4",x"49"),
   599 => (x"aa",x"71",x"41",x"20"),
   600 => (x"26",x"87",x"f9",x"05"),
   601 => (x"fe",x"f9",x"c2",x"4a"),
   602 => (x"87",x"eb",x"f6",x"49"),
   603 => (x"c4",x"05",x"98",x"70"),
   604 => (x"d4",x"e6",x"c2",x"87"),
   605 => (x"fe",x"49",x"c0",x"4b"),
   606 => (x"73",x"87",x"e5",x"c5"),
   607 => (x"87",x"c7",x"fe",x"48"),
   608 => (x"00",x"20",x"20",x"20"),
   609 => (x"45",x"54",x"4f",x"4a"),
   610 => (x"20",x"20",x"4f",x"47"),
   611 => (x"00",x"20",x"20",x"20"),
   612 => (x"00",x"43",x"52",x"41"),
   613 => (x"20",x"43",x"52",x"41"),
   614 => (x"20",x"74",x"6f",x"6e"),
   615 => (x"6e",x"75",x"6f",x"66"),
   616 => (x"4c",x"20",x"2e",x"64"),
   617 => (x"20",x"64",x"61",x"6f"),
   618 => (x"00",x"43",x"52",x"41"),
   619 => (x"87",x"e8",x"eb",x"1e"),
   620 => (x"f8",x"87",x"ef",x"fb"),
   621 => (x"16",x"4f",x"26",x"87"),
   622 => (x"2e",x"25",x"26",x"1e"),
   623 => (x"2e",x"3e",x"3d",x"36"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

