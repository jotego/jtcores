/*  This file is part of JTFRAME.
    JTFRAME program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTFRAME program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTFRAME.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 8-5-2021 */

// ctrl+shift selects sys info
// alt+shift selects target info

module jtframe_debug #(
    parameter COLORW=4
) (
    input              clk,
    input              rst,

    input              shift,         // count step 16, instead of 1
    input              ctrl,          // reset debug_bus
    input              alt,
    input              toggle_view,
    input        [1:0] debug_plus,
    input        [1:0] debug_minus,
    input        [7:0] key_digit,
    // overlay the value on video
    input              pxl_cen,
    input [COLORW-1:0] rin,
    input [COLORW-1:0] gin,
    input [COLORW-1:0] bin,
    input              lhbl,
    input              lvbl,
    input              dip_flip,

    // combinational output
    output [COLORW-1:0] rout,
    output [COLORW-1:0] gout,
    output [COLORW-1:0] bout,
    // debug features
    output        [7:0] debug_bus,
    input         [7:0] debug_view, // an 8-bit signal that will be shown over the game image
    input         [7:0] sys_info,   // system information generated within JTFRAME, not the game
    input         [7:0] target_info,  // system information generated by the JTFRAME target, not the game
    input         [7:0] snd_vol,
    input               snd_mode
);

wire [2:0] color;
wire [7:0] view_bin, view_hex, msg;
wire [8:0] h, v;
wire [1:0] view_mode;
wire       split_binhex, hex_en, bin_en;

jtframe_debug_ctrl u_ctrl(
    .clk        ( clk           ),
    .pxl_cen    ( pxl_cen       ),

    .debug_bus  ( debug_bus     ),
    .view_bin   ( view_bin      ),
    .view_hex   ( view_hex      ),
    .v          ( v             ),
    .h          ( h             ),
    .view_mode  ( view_mode     ),

    .split_binhex(split_binhex  ),

    .hex_en     ( hex_en        ),
    .bin_en     ( bin_en        ),
    .color      ( color         ),
    .msg        ( msg           )
);

jtframe_debug_viewmux u_viewmux(
    .rst        ( rst           ),
    .clk        ( clk           ),
    .toggle     ( toggle_view   ),

    .debug_view ( debug_view    ),
    .sys_info   ( sys_info      ),
    .target_info( target_info   ),

    .snd_mode    ( snd_mode     ),
    .snd_vol     ( snd_vol      ),
    .split_binhex(split_binhex  ),

    .view_bin   ( view_bin      ),
    .view_hex   ( view_hex      ),
    .sel        ( view_mode     )
);

jtframe_binhex_overlay #(.COLORW(COLORW)) u_overlay(
    .clk        ( clk         ),
    .v          ( v           ),
    .h          ( h           ),

    .bin_en     ( bin_en      ),
    .hex_en     ( hex_en      ),
    .din        ( msg         ),
    .color      ( color       ),

    .rin        ( rin         ),
    .gin        ( gin         ),
    .bin        ( bin         ),

    .rout       ( rout        ),
    .gout       ( gout        ),
    .bout       ( bout        )
);

jtframe_video_counter u_vcounters(
    .rst        ( rst         ),
    .clk        ( clk         ),
    .pxl_cen    ( pxl_cen     ),

    .lhbl       ( lhbl        ),
    .lvbl       ( lvbl        ),
    .hs         ( 1'b0        ), // not needed if len outputs are not used
    .vs         ( 1'b0        ), // not needed if len outputs are not used
    .flip       ( dip_flip    ),

    .v          ( v           ),
    .h          ( h           ),

    .hbs_len    (             ),
    .hsy_len    (             ),
    .hsa_len    (             ),

    .vbs_len    (             ),
    .vsy_len    (             ),
    .vsa_len    (             ),
    .rdy        (             )
);

jtframe_debug_bus u_debug_bus(
    .rst        ( rst         ),
    .clk        ( clk         ),
    .shift      ( shift       ),
    .ctrl       ( ctrl        ),
    .inc        ( debug_plus  ),
    .dec        ( debug_minus ),
    .key_digit  ( key_digit   ),
    .debug_bus  ( debug_bus   )
);

endmodule