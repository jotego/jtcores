-------------------------------------------------------------------------------
--
-- The UPI-41 BUS unit.
-- Implements the BUS port logic.
--
-- Copyright (c) 2004-2022, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration upi41_db_bus_rtl_c0 of upi41_db_bus is

  for rtl
  end for;

end upi41_db_bus_rtl_c0;
