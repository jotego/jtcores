../../cps1/hdl/turbo.vh