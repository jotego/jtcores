localparam [2:0] XMEN=3'd2;