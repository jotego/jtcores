/*  This file is part of JTFRAME.
    JTFRAME program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTFRAME program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTFRAME.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 26-1-2025 */

module jtframe_debug_viewmux(
    input            clk,
    input            toggle,

    input      [7:0] debug_view, // an 8-bit signal that will be shown over the game image
    input      [7:0] sys_info,   // system information generated within JTFRAME, not the game
    input      [7:0] target_info,  // system information generated by the JTFRAME target, not the game
    input            snd_mode,
    input      [7:0] snd_vol,

    output reg       split_binhex=0,
    output reg [1:0] sel=0,
    output reg [7:0] view_bin=0,
    output reg [7:0] view_hex=0
);    

`include "jtframe_debug.vh"

reg  [7:0] mux;
reg        toggle_l;

always @(posedge clk) begin
    toggle_l <= toggle;

    if( toggle && !toggle_l ) begin
        sel <= sel==2 ? 2'd0 : sel+1'd1;
    end
end

always @(posedge clk) begin
    case( sel )
        default:     mux <= debug_view;
        SYS_INFO:    mux <= sys_info;
        TARGET_INFO: mux <= target_info;
    endcase
    split_binhex <= sel==SYS_INFO && snd_mode;

    view_bin <= mux;
    view_hex <= split_binhex ? snd_vol : view_bin;
end

endmodule