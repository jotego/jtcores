`timescale 1ns/1ps

module test;

reg clk, rst;

initial begin
    clk=0;
    forever #83.33 clk = ~clk;
end

integer hcnt=0,vcnt=0, frame=0;

wire lhbl = ~(hcnt>=160 && hcnt<180);
wire lvbl = ~(vcnt>=152 && vcnt<160);

always @(posedge clk) begin
    hcnt <= hcnt==180 ? 0 : hcnt+1;
    if( hcnt==170 ) begin
        vcnt <= vcnt==160 ? 0 : vcnt+1;
        if( vcnt==158 ) frame<=frame+1;
        if( frame==3 ) $finish;
    end
end

initial begin
    $dumpfile("test.lxt");
    $dumpvars;
    $dumpon;
end

initial begin
    rst=0;
    hcnt=0;
    vcnt=0;
    frame=0;
    #10 rst=1;
    #500 rst=0;
    #110000000 $finish;
end

jtframe_debug uut(
    .clk        ( clk   ),
    .rst        ( rst   ),

    .shift      ( 0     ),         // count step 16, instead of 1
    .ctrl       ( 0     ),          // reset debug_bus
    .alt        ( 0     ),
    .debug_plus ( 1'b1  ),
    .debug_minus( 0     ),
    .debug_rst  ( 0     ),
    .key_gfx    ( 0     ),
    .key_digit  ( 0     ),
    // overlay the value on video
    .pxl_cen    ( 1     ),
    .rin        ( 0     ),
    .gin        ( 0     ),
    .bin        ( 0     ),
    .lhbl       ( lhbl  ),
    .lvbl       ( lvbl  ),
    .dip_flip   ( 0     ),

    // combinational output
    .rout       (       ),
    .gout       (       ),
    .bout       (       ),
    // debug features
    .debug_bus  (       ),
    .debug_view ( 8'h10 ), // an 8-bit signal that will be shown over the game image
    .sys_info   ( 0     ),   // system information generated within JTFRAME, not the game
    .target_info( 0     ),  // system information generated by the JTFRAME target, not the game
    .gfx_en     (       )
);

endmodule