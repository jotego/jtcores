/*  This file is part of JTCORES1.
    JTCORES1 program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTCORES1.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 16-2-2021 */


module jtcps2_sbox_fn1_r1(
    input  [ 7:0] din,
    input  [23:0] key,
    output [ 7:0] dout
);

    jtcps2_sbox #(
        .LUT( {
        2'd3, 2'd1, 2'd0, 2'd2, 2'd3, 2'd1, 2'd3, 2'd2, 
        2'd2, 2'd2, 2'd3, 2'd2, 2'd1, 2'd2, 2'd2, 2'd1, 
        2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd3, 2'd1, 2'd1, 
        2'd1, 2'd3, 2'd1, 2'd3, 2'd0, 2'd0, 2'd2, 2'd2, 
        2'd2, 2'd1, 2'd1, 2'd1, 2'd2, 2'd3, 2'd3, 2'd2, 
        2'd2, 2'd2, 2'd3, 2'd1, 2'd2, 2'd1, 2'd1, 2'd1, 
        2'd2, 2'd1, 2'd3, 2'd0, 2'd3, 2'd0, 2'd2, 2'd3, 
        2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd2, 2'd2, 2'd0
        } ),
        .LOC( { 3'd0, 3'd0, 3'd6, 3'd5, 3'd4, 3'd3 } ),
        .OK ( 6'b00_1111 ))
    u_sbox_fn1_r1_0(
        .din ( din                  ),
        .key ( key[ 5:0 ]           ),
        .dout( { dout[6], dout[3] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd0, 2'd3, 2'd2, 2'd3, 2'd1, 2'd3, 2'd2, 
        2'd2, 2'd2, 2'd3, 2'd1, 2'd1, 2'd3, 2'd2, 2'd3, 
        2'd1, 2'd2, 2'd1, 2'd0, 2'd2, 2'd1, 2'd1, 2'd1, 
        2'd1, 2'd3, 2'd3, 2'd3, 2'd2, 2'd3, 2'd1, 2'd0, 
        2'd3, 2'd3, 2'd3, 2'd0, 2'd3, 2'd2, 2'd2, 2'd1, 
        2'd2, 2'd0, 2'd0, 2'd0, 2'd3, 2'd1, 2'd3, 2'd2, 
        2'd3, 2'd2, 2'd0, 2'd0, 2'd0, 2'd1, 2'd2, 2'd1, 
        2'd1, 2'd1, 2'd1, 2'd2, 2'd2, 2'd2, 2'd0, 2'd3
        } ),
        .LOC( { 3'd0, 3'd7, 3'd4, 3'd2, 3'd1, 3'd0 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn1_r1_1(
        .din ( din                  ),
        .key ( key[11:6 ]           ),
        .dout( { dout[7], dout[2] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd0, 2'd0, 2'd2, 2'd2, 2'd0, 2'd2, 2'd1, 
        2'd1, 2'd1, 2'd3, 2'd1, 2'd3, 2'd2, 2'd1, 2'd3, 
        2'd0, 2'd1, 2'd2, 2'd0, 2'd1, 2'd0, 2'd1, 2'd2, 
        2'd0, 2'd2, 2'd0, 2'd1, 2'd2, 2'd1, 2'd3, 2'd2, 
        2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd2, 2'd0, 
        2'd2, 2'd0, 2'd3, 2'd2, 2'd1, 2'd0, 2'd1, 2'd0, 
        2'd3, 2'd2, 2'd3, 2'd3, 2'd0, 2'd2, 2'd1, 2'd3, 
        2'd2, 2'd2, 2'd0, 2'd1, 2'd1, 2'd3, 2'd0, 2'd3
        } ),
        .LOC( { 3'd7, 3'd6, 3'd3, 3'd2, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r1_2(
        .din ( din                  ),
        .key ( key[17:12]           ),
        .dout( { dout[1], dout[0] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd3, 2'd3, 2'd1, 2'd1, 2'd0, 2'd3, 2'd0, 2'd0, 
        2'd3, 2'd3, 2'd1, 2'd2, 2'd0, 2'd2, 2'd3, 2'd3, 
        2'd0, 2'd2, 2'd3, 2'd2, 2'd2, 2'd1, 2'd1, 2'd3, 
        2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd2, 
        2'd2, 2'd0, 2'd0, 2'd0, 2'd3, 2'd1, 2'd0, 2'd1, 
        2'd0, 2'd1, 2'd2, 2'd3, 2'd3, 2'd1, 2'd2, 2'd2, 
        2'd1, 2'd2, 2'd3, 2'd1, 2'd2, 2'd3, 2'd2, 2'd1, 
        2'd1, 2'd2, 2'd2, 2'd0, 2'd3, 2'd0, 2'd2, 2'd3
        } ),
        .LOC( { 3'd7, 3'd6, 3'd5, 3'd3, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r1_3(
        .din ( din                  ),
        .key ( key[23:18]           ),
        .dout( { dout[5], dout[4] } )
    );

endmodule


module jtcps2_sbox_fn1_r2(
    input  [ 7:0] din,
    input  [23:0] key,
    output [ 7:0] dout
);

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd3, 2'd1, 2'd0, 2'd2, 2'd1, 2'd2, 2'd1, 
        2'd2, 2'd2, 2'd1, 2'd0, 2'd3, 2'd1, 2'd0, 2'd3, 
        2'd2, 2'd1, 2'd2, 2'd3, 2'd1, 2'd0, 2'd3, 2'd3, 
        2'd0, 2'd2, 2'd1, 2'd0, 2'd1, 2'd2, 2'd2, 2'd0, 
        2'd2, 2'd1, 2'd3, 2'd2, 2'd2, 2'd3, 2'd2, 2'd3, 
        2'd3, 2'd3, 2'd1, 2'd3, 2'd3, 2'd0, 2'd3, 2'd1, 
        2'd3, 2'd1, 2'd2, 2'd0, 2'd1, 2'd0, 2'd3, 2'd0, 
        2'd1, 2'd3, 2'd0, 2'd3, 2'd0, 2'd2, 2'd3, 2'd3
        } ),
        .LOC( { 3'd0, 3'd6, 3'd3, 3'd2, 3'd1, 3'd0 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn1_r2_0(
        .din ( din                  ),
        .key ( key[ 5:0 ]           ),
        .dout( { dout[6], dout[1] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd2, 2'd0, 2'd3, 2'd2, 2'd3, 2'd0, 2'd2, 
        2'd3, 2'd1, 2'd2, 2'd1, 2'd3, 2'd2, 2'd1, 2'd0, 
        2'd3, 2'd0, 2'd1, 2'd2, 2'd1, 2'd2, 2'd1, 2'd2, 
        2'd3, 2'd2, 2'd0, 2'd1, 2'd0, 2'd2, 2'd2, 2'd2, 
        2'd3, 2'd1, 2'd2, 2'd3, 2'd2, 2'd1, 2'd0, 2'd1, 
        2'd0, 2'd1, 2'd2, 2'd2, 2'd1, 2'd0, 2'd3, 2'd3, 
        2'd2, 2'd3, 2'd2, 2'd0, 2'd0, 2'd2, 2'd0, 2'd1, 
        2'd1, 2'd0, 2'd3, 2'd1, 2'd2, 2'd3, 2'd2, 2'd1
        } ),
        .LOC( { 3'd0, 3'd7, 3'd6, 3'd5, 3'd4, 3'd2 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn1_r2_1(
        .din ( din                  ),
        .key ( key[11:6 ]           ),
        .dout( { dout[7], dout[5] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd3, 2'd1, 2'd3, 2'd2, 2'd3, 2'd0, 2'd0, 2'd2, 
        2'd2, 2'd1, 2'd1, 2'd1, 2'd2, 2'd2, 2'd2, 2'd1, 
        2'd0, 2'd0, 2'd1, 2'd1, 2'd2, 2'd3, 2'd3, 2'd1, 
        2'd0, 2'd3, 2'd1, 2'd3, 2'd0, 2'd3, 2'd1, 2'd1, 
        2'd2, 2'd2, 2'd2, 2'd3, 2'd3, 2'd3, 2'd0, 2'd1, 
        2'd3, 2'd2, 2'd2, 2'd2, 2'd1, 2'd3, 2'd1, 2'd1, 
        2'd0, 2'd0, 2'd3, 2'd1, 2'd2, 2'd2, 2'd2, 2'd0, 
        2'd1, 2'd0, 2'd1, 2'd1, 2'd2, 2'd0, 2'd1, 2'd0
        } ),
        .LOC( { 3'd7, 3'd5, 3'd4, 3'd3, 3'd2, 3'd1 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r2_2(
        .din ( din                  ),
        .key ( key[17:12]           ),
        .dout( { dout[3], dout[0] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd3, 2'd3, 2'd2, 2'd1, 2'd0, 2'd1, 2'd3, 2'd1, 
        2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd0, 
        2'd3, 2'd1, 2'd1, 2'd2, 2'd2, 2'd2, 2'd1, 2'd2, 
        2'd0, 2'd2, 2'd3, 2'd0, 2'd3, 2'd3, 2'd3, 2'd1, 
        2'd0, 2'd3, 2'd0, 2'd3, 2'd0, 2'd3, 2'd0, 2'd0, 
        2'd0, 2'd1, 2'd2, 2'd1, 2'd0, 2'd3, 2'd3, 2'd1, 
        2'd1, 2'd3, 2'd0, 2'd1, 2'd1, 2'd1, 2'd2, 2'd1, 
        2'd0, 2'd2, 2'd3, 2'd3, 2'd3, 2'd0, 2'd1, 2'd2
        } ),
        .LOC( { 3'd7, 3'd6, 3'd4, 3'd3, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r2_3(
        .din ( din                  ),
        .key ( key[23:18]           ),
        .dout( { dout[4], dout[2] } )
    );

endmodule


module jtcps2_sbox_fn1_r3(
    input  [ 7:0] din,
    input  [23:0] key,
    output [ 7:0] dout
);

    jtcps2_sbox #(
        .LUT( {
        2'd3, 2'd3, 2'd3, 2'd3, 2'd3, 2'd1, 2'd3, 2'd0, 
        2'd0, 2'd0, 2'd2, 2'd0, 2'd1, 2'd0, 2'd0, 2'd2, 
        2'd3, 2'd3, 2'd1, 2'd0, 2'd2, 2'd3, 2'd1, 2'd0, 
        2'd3, 2'd3, 2'd2, 2'd1, 2'd1, 2'd0, 2'd0, 2'd3, 
        2'd3, 2'd2, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd3, 
        2'd0, 2'd1, 2'd2, 2'd2, 2'd3, 2'd2, 2'd1, 2'd0, 
        2'd2, 2'd3, 2'd0, 2'd0, 2'd0, 2'd2, 2'd0, 2'd2, 
        2'd0, 2'd1, 2'd1, 2'd3, 2'd3, 2'd0, 2'd0, 2'd0
        } ),
        .LOC( { 3'd0, 3'd7, 3'd6, 3'd5, 3'd1, 3'd0 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn1_r3_0(
        .din ( din                  ),
        .key ( key[ 5:0 ]           ),
        .dout( { dout[5], dout[0] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd3, 2'd1, 2'd1, 2'd1, 2'd2, 2'd0, 2'd3, 2'd1, 
        2'd3, 2'd1, 2'd2, 2'd0, 2'd3, 2'd2, 2'd2, 2'd1, 
        2'd0, 2'd1, 2'd2, 2'd0, 2'd1, 2'd3, 2'd2, 2'd3, 
        2'd0, 2'd3, 2'd3, 2'd2, 2'd1, 2'd2, 2'd0, 2'd3, 
        2'd1, 2'd2, 2'd2, 2'd1, 2'd2, 2'd0, 2'd1, 2'd0, 
        2'd0, 2'd1, 2'd1, 2'd1, 2'd3, 2'd2, 2'd0, 2'd1, 
        2'd2, 2'd0, 2'd2, 2'd3, 2'd0, 2'd3, 2'd2, 2'd2, 
        2'd0, 2'd3, 2'd2, 2'd0, 2'd3, 2'd2, 2'd3, 2'd2
        } ),
        .LOC( { 3'd0, 3'd7, 3'd6, 3'd4, 3'd3, 3'd2 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn1_r3_1(
        .din ( din                  ),
        .key ( key[11:6 ]           ),
        .dout( { dout[7], dout[6] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd0, 2'd0, 2'd2, 2'd3, 2'd0, 2'd0, 2'd0, 
        2'd0, 2'd3, 2'd2, 2'd0, 2'd0, 2'd1, 2'd1, 2'd3, 
        2'd0, 2'd3, 2'd1, 2'd0, 2'd2, 2'd1, 2'd1, 2'd3, 
        2'd2, 2'd1, 2'd0, 2'd0, 2'd2, 2'd1, 2'd1, 2'd2, 
        2'd0, 2'd3, 2'd0, 2'd0, 2'd0, 2'd2, 2'd1, 2'd3, 
        2'd2, 2'd0, 2'd0, 2'd2, 2'd0, 2'd1, 2'd3, 2'd2, 
        2'd1, 2'd0, 2'd0, 2'd2, 2'd2, 2'd2, 2'd1, 2'd2, 
        2'd2, 2'd1, 2'd3, 2'd1, 2'd1, 2'd2, 2'd0, 2'd3
        } ),
        .LOC( { 3'd6, 3'd5, 3'd4, 3'd3, 3'd2, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r3_2(
        .din ( din                  ),
        .key ( key[17:12]           ),
        .dout( { dout[4], dout[1] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd1, 2'd1, 2'd3, 2'd0, 2'd3, 2'd2, 2'd0, 
        2'd1, 2'd3, 2'd2, 2'd2, 2'd3, 2'd3, 2'd3, 2'd0, 
        2'd0, 2'd1, 2'd2, 2'd2, 2'd2, 2'd3, 2'd2, 2'd1, 
        2'd1, 2'd2, 2'd0, 2'd3, 2'd0, 2'd3, 2'd3, 2'd1, 
        2'd2, 2'd3, 2'd3, 2'd0, 2'd1, 2'd2, 2'd2, 2'd0, 
        2'd0, 2'd1, 2'd1, 2'd3, 2'd3, 2'd0, 2'd1, 2'd1, 
        2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd2, 2'd3, 2'd3, 
        2'd2, 2'd3, 2'd1, 2'd2, 2'd0, 2'd0, 2'd1, 2'd0
        } ),
        .LOC( { 3'd7, 3'd5, 3'd3, 3'd2, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r3_3(
        .din ( din                  ),
        .key ( key[23:18]           ),
        .dout( { dout[3], dout[2] } )
    );

endmodule


module jtcps2_sbox_fn1_r4(
    input  [ 7:0] din,
    input  [23:0] key,
    output [ 7:0] dout
);

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd3, 2'd3, 2'd1, 2'd0, 2'd3, 2'd1, 2'd3, 
        2'd0, 2'd3, 2'd1, 2'd2, 2'd0, 2'd0, 2'd0, 2'd2, 
        2'd2, 2'd1, 2'd0, 2'd2, 2'd3, 2'd2, 2'd1, 2'd3, 
        2'd2, 2'd3, 2'd1, 2'd2, 2'd3, 2'd0, 2'd1, 2'd0, 
        2'd2, 2'd1, 2'd0, 2'd2, 2'd3, 2'd2, 2'd3, 2'd0, 
        2'd3, 2'd2, 2'd1, 2'd2, 2'd1, 2'd0, 2'd3, 2'd3, 
        2'd2, 2'd0, 2'd2, 2'd1, 2'd0, 2'd3, 2'd2, 2'd3, 
        2'd3, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1
        } ),
        .LOC( { 3'd7, 3'd5, 3'd4, 3'd3, 3'd2, 3'd1 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r4_0(
        .din ( din                  ),
        .key ( key[ 5:0 ]           ),
        .dout( { dout[4], dout[0] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd1, 2'd2, 2'd2, 2'd3, 2'd3, 2'd1, 2'd0, 
        2'd0, 2'd1, 2'd1, 2'd3, 2'd1, 2'd0, 2'd3, 2'd0, 
        2'd1, 2'd0, 2'd2, 2'd0, 2'd2, 2'd0, 2'd3, 2'd0, 
        2'd3, 2'd0, 2'd3, 2'd2, 2'd0, 2'd3, 2'd1, 2'd1, 
        2'd0, 2'd0, 2'd3, 2'd3, 2'd2, 2'd2, 2'd0, 2'd1, 
        2'd0, 2'd2, 2'd0, 2'd0, 2'd1, 2'd3, 2'd2, 2'd2, 
        2'd2, 2'd1, 2'd3, 2'd0, 2'd3, 2'd1, 2'd3, 2'd3, 
        2'd2, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0, 2'd0, 2'd3
        } ),
        .LOC( { 3'd6, 3'd5, 3'd3, 3'd2, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r4_1(
        .din ( din                  ),
        .key ( key[11:6 ]           ),
        .dout( { dout[3], dout[1] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd3, 2'd1, 2'd1, 2'd3, 2'd3, 2'd2, 2'd1, 
        2'd3, 2'd0, 2'd3, 2'd2, 2'd1, 2'd1, 2'd1, 2'd2, 
        2'd1, 2'd0, 2'd0, 2'd2, 2'd2, 2'd0, 2'd1, 2'd1, 
        2'd2, 2'd2, 2'd2, 2'd0, 2'd3, 2'd2, 2'd0, 2'd3, 
        2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd2, 2'd3, 
        2'd2, 2'd3, 2'd3, 2'd2, 2'd2, 2'd1, 2'd0, 2'd3, 
        2'd0, 2'd3, 2'd0, 2'd0, 2'd2, 2'd3, 2'd0, 2'd2, 
        2'd1, 2'd3, 2'd1, 2'd0, 2'd2, 2'd1, 2'd1, 2'd0
        } ),
        .LOC( { 3'd7, 3'd6, 3'd5, 3'd4, 3'd2, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r4_2(
        .din ( din                  ),
        .key ( key[17:12]           ),
        .dout( { dout[6], dout[2] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd0, 2'd3, 2'd2, 2'd1, 2'd2, 2'd2, 2'd2, 
        2'd0, 2'd0, 2'd0, 2'd3, 2'd0, 2'd0, 2'd1, 2'd3, 
        2'd0, 2'd3, 2'd2, 2'd3, 2'd2, 2'd3, 2'd3, 2'd0, 
        2'd1, 2'd1, 2'd2, 2'd1, 2'd3, 2'd1, 2'd1, 2'd1, 
        2'd3, 2'd3, 2'd1, 2'd2, 2'd0, 2'd0, 2'd2, 2'd3, 
        2'd3, 2'd2, 2'd2, 2'd0, 2'd3, 2'd3, 2'd1, 2'd0, 
        2'd2, 2'd0, 2'd2, 2'd3, 2'd1, 2'd1, 2'd2, 2'd2, 
        2'd3, 2'd0, 2'd1, 2'd0, 2'd2, 2'd2, 2'd1, 2'd0
        } ),
        .LOC( { 3'd7, 3'd6, 3'd4, 3'd3, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn1_r4_3(
        .din ( din                  ),
        .key ( key[23:18]           ),
        .dout( { dout[7], dout[5] } )
    );

endmodule


module jtcps2_sbox_fn2_r1(
    input  [ 7:0] din,
    input  [23:0] key,
    output [ 7:0] dout
);

    jtcps2_sbox #(
        .LUT( {
        2'd1, 2'd3, 2'd1, 2'd1, 2'd3, 2'd1, 2'd2, 2'd2, 
        2'd1, 2'd1, 2'd3, 2'd0, 2'd2, 2'd0, 2'd1, 2'd1, 
        2'd2, 2'd1, 2'd0, 2'd3, 2'd2, 2'd0, 2'd3, 2'd0, 
        2'd3, 2'd3, 2'd2, 2'd2, 2'd1, 2'd0, 2'd1, 2'd0, 
        2'd0, 2'd3, 2'd1, 2'd2, 2'd0, 2'd3, 2'd2, 2'd2, 
        2'd2, 2'd0, 2'd2, 2'd0, 2'd2, 2'd1, 2'd0, 2'd2, 
        2'd1, 2'd0, 2'd2, 2'd3, 2'd1, 2'd0, 2'd1, 2'd1, 
        2'd3, 2'd0, 2'd0, 2'd3, 2'd0, 2'd2, 2'd0, 2'd2
        } ),
        .LOC( { 3'd0, 3'd7, 3'd5, 3'd4, 3'd3, 3'd0 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn2_r1_0(
        .din ( din                  ),
        .key ( key[ 5:0 ]           ),
        .dout( { dout[7], dout[6] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd3, 2'd1, 2'd1, 2'd1, 2'd3, 2'd2, 2'd2, 
        2'd3, 2'd3, 2'd3, 2'd0, 2'd2, 2'd1, 2'd1, 2'd3, 
        2'd2, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd2, 2'd2, 
        2'd2, 2'd2, 2'd2, 2'd2, 2'd3, 2'd1, 2'd3, 2'd1, 
        2'd1, 2'd1, 2'd3, 2'd3, 2'd3, 2'd1, 2'd0, 2'd2, 
        2'd2, 2'd2, 2'd2, 2'd0, 2'd2, 2'd2, 2'd3, 2'd1, 
        2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd2, 2'd0, 2'd3, 
        2'd1, 2'd0, 2'd2, 2'd0, 2'd3, 2'd0, 2'd1, 2'd1
        } ),
        .LOC( { 3'd0, 3'd6, 3'd4, 3'd3, 3'd2, 3'd1 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn2_r1_1(
        .din ( din                  ),
        .key ( key[11:6 ]           ),
        .dout( { dout[5], dout[3] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd3, 2'd1, 2'd1, 2'd3, 2'd1, 2'd2, 2'd3, 2'd1, 
        2'd0, 2'd2, 2'd3, 2'd2, 2'd0, 2'd0, 2'd0, 2'd3, 
        2'd1, 2'd0, 2'd3, 2'd2, 2'd3, 2'd2, 2'd0, 2'd0, 
        2'd0, 2'd2, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd2, 
        2'd2, 2'd0, 2'd0, 2'd0, 2'd2, 2'd1, 2'd3, 2'd2, 
        2'd1, 2'd0, 2'd0, 2'd2, 2'd1, 2'd3, 2'd2, 2'd1, 
        2'd1, 2'd2, 2'd1, 2'd0, 2'd1, 2'd2, 2'd2, 2'd1, 
        2'd3, 2'd3, 2'd3, 2'd3, 2'd2, 2'd2, 2'd0, 2'd1
        } ),
        .LOC( { 3'd7, 3'd6, 3'd5, 3'd4, 3'd2, 3'd1 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r1_2(
        .din ( din                  ),
        .key ( key[17:12]           ),
        .dout( { dout[4], dout[1] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd2, 2'd2, 2'd3, 2'd1, 2'd0, 2'd3, 2'd0, 
        2'd0, 2'd0, 2'd3, 2'd1, 2'd2, 2'd1, 2'd3, 2'd3, 
        2'd2, 2'd2, 2'd2, 2'd0, 2'd1, 2'd0, 2'd0, 2'd3, 
        2'd1, 2'd2, 2'd1, 2'd0, 2'd0, 2'd0, 2'd3, 2'd2, 
        2'd1, 2'd0, 2'd3, 2'd3, 2'd0, 2'd0, 2'd0, 2'd3, 
        2'd2, 2'd0, 2'd0, 2'd1, 2'd3, 2'd0, 2'd3, 2'd2, 
        2'd1, 2'd2, 2'd3, 2'd3, 2'd1, 2'd1, 2'd2, 2'd3, 
        2'd1, 2'd3, 2'd2, 2'd3, 2'd0, 2'd3, 2'd3, 2'd1
        } ),
        .LOC( { 3'd7, 3'd6, 3'd5, 3'd3, 3'd2, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r1_3(
        .din ( din                  ),
        .key ( key[23:18]           ),
        .dout( { dout[2], dout[0] } )
    );

endmodule


module jtcps2_sbox_fn2_r2(
    input  [ 7:0] din,
    input  [23:0] key,
    output [ 7:0] dout
);

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd1, 2'd1, 2'd2, 2'd1, 2'd2, 2'd1, 2'd1, 
        2'd0, 2'd0, 2'd2, 2'd0, 2'd0, 2'd3, 2'd3, 2'd0, 
        2'd2, 2'd0, 2'd1, 2'd1, 2'd1, 2'd2, 2'd1, 2'd3, 
        2'd0, 2'd3, 2'd3, 2'd1, 2'd1, 2'd2, 2'd2, 2'd2, 
        2'd3, 2'd2, 2'd0, 2'd2, 2'd2, 2'd2, 2'd1, 2'd3, 
        2'd3, 2'd2, 2'd3, 2'd2, 2'd1, 2'd0, 2'd1, 2'd1, 
        2'd3, 2'd0, 2'd3, 2'd1, 2'd1, 2'd0, 2'd0, 2'd3, 
        2'd1, 2'd3, 2'd0, 2'd3, 2'd0, 2'd3, 2'd1, 2'd3
        } ),
        .LOC( { 3'd0, 3'd0, 3'd6, 3'd4, 3'd2, 3'd0 } ),
        .OK ( 6'b00_1111 ))
    u_sbox_fn2_r2_0(
        .din ( din                  ),
        .key ( key[ 5:0 ]           ),
        .dout( { dout[6], dout[4] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd2, 2'd1, 2'd0, 2'd0, 2'd3, 2'd1, 2'd1, 
        2'd3, 2'd0, 2'd3, 2'd3, 2'd2, 2'd0, 2'd1, 2'd3, 
        2'd3, 2'd2, 2'd0, 2'd2, 2'd1, 2'd2, 2'd0, 2'd2, 
        2'd1, 2'd1, 2'd0, 2'd2, 2'd1, 2'd0, 2'd3, 2'd2, 
        2'd0, 2'd1, 2'd0, 2'd2, 2'd2, 2'd1, 2'd2, 2'd3, 
        2'd3, 2'd3, 2'd1, 2'd2, 2'd2, 2'd1, 2'd3, 2'd0, 
        2'd3, 2'd2, 2'd0, 2'd2, 2'd1, 2'd1, 2'd1, 2'd3, 
        2'd2, 2'd1, 2'd2, 2'd3, 2'd3, 2'd0, 2'd3, 2'd0
        } ),
        .LOC( { 3'd7, 3'd6, 3'd5, 3'd4, 3'd3, 3'd1 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r2_1(
        .din ( din                  ),
        .key ( key[11:6 ]           ),
        .dout( { dout[3], dout[0] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd1, 2'd2, 2'd0, 2'd1, 2'd2, 2'd3, 2'd2, 2'd1, 
        2'd2, 2'd2, 2'd0, 2'd2, 2'd2, 2'd3, 2'd0, 2'd3, 
        2'd3, 2'd0, 2'd3, 2'd2, 2'd1, 2'd0, 2'd2, 2'd1, 
        2'd1, 2'd1, 2'd0, 2'd1, 2'd2, 2'd2, 2'd3, 2'd3, 
        2'd1, 2'd3, 2'd2, 2'd1, 2'd1, 2'd0, 2'd0, 2'd3, 
        2'd0, 2'd1, 2'd1, 2'd2, 2'd3, 2'd2, 2'd2, 2'd1, 
        2'd3, 2'd0, 2'd1, 2'd1, 2'd2, 2'd2, 2'd2, 2'd1, 
        2'd0, 2'd1, 2'd2, 2'd3, 2'd1, 2'd2, 2'd0, 2'd0
        } ),
        .LOC( { 3'd7, 3'd5, 3'd4, 3'd3, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r2_2(
        .din ( din                  ),
        .key ( key[17:12]           ),
        .dout( { dout[7], dout[1] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd2, 2'd3, 2'd2, 2'd2, 2'd1, 2'd0, 2'd0, 
        2'd3, 2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 
        2'd1, 2'd3, 2'd2, 2'd3, 2'd0, 2'd2, 2'd3, 2'd0, 
        2'd0, 2'd0, 2'd1, 2'd1, 2'd3, 2'd3, 2'd3, 2'd2, 
        2'd2, 2'd1, 2'd2, 2'd2, 2'd0, 2'd0, 2'd2, 2'd2, 
        2'd1, 2'd3, 2'd2, 2'd1, 2'd3, 2'd2, 2'd3, 2'd3, 
        2'd0, 2'd3, 2'd2, 2'd3, 2'd0, 2'd2, 2'd3, 2'd1, 
        2'd0, 2'd2, 2'd2, 2'd0, 2'd2, 2'd1, 2'd2, 2'd0
        } ),
        .LOC( { 3'd7, 3'd6, 3'd5, 3'd3, 3'd2, 3'd1 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r2_3(
        .din ( din                  ),
        .key ( key[23:18]           ),
        .dout( { dout[5], dout[2] } )
    );

endmodule


module jtcps2_sbox_fn2_r3(
    input  [ 7:0] din,
    input  [23:0] key,
    output [ 7:0] dout
);

    jtcps2_sbox #(
        .LUT( {
        2'd1, 2'd3, 2'd3, 2'd2, 2'd0, 2'd1, 2'd2, 2'd1, 
        2'd0, 2'd3, 2'd3, 2'd3, 2'd0, 2'd0, 2'd0, 2'd0, 
        2'd0, 2'd2, 2'd3, 2'd3, 2'd3, 2'd2, 2'd2, 2'd0, 
        2'd2, 2'd2, 2'd3, 2'd1, 2'd1, 2'd2, 2'd1, 2'd1, 
        2'd2, 2'd1, 2'd2, 2'd3, 2'd2, 2'd0, 2'd1, 2'd1, 
        2'd0, 2'd0, 2'd1, 2'd3, 2'd3, 2'd0, 2'd2, 2'd0, 
        2'd1, 2'd0, 2'd0, 2'd3, 2'd3, 2'd1, 2'd2, 2'd2, 
        2'd3, 2'd1, 2'd3, 2'd2, 2'd1, 2'd2, 2'd1, 2'd2
        } ),
        .LOC( { 3'd0, 3'd0, 3'd6, 3'd4, 3'd3, 3'd2 } ),
        .OK ( 6'b00_1111 ))
    u_sbox_fn2_r3_0(
        .din ( din                  ),
        .key ( key[ 5:0 ]           ),
        .dout( { dout[5], dout[3] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd0, 2'd3, 2'd2, 2'd2, 2'd2, 2'd0, 2'd1, 
        2'd3, 2'd3, 2'd0, 2'd2, 2'd3, 2'd1, 2'd3, 2'd1, 
        2'd0, 2'd0, 2'd2, 2'd0, 2'd0, 2'd1, 2'd0, 2'd2, 
        2'd2, 2'd0, 2'd0, 2'd1, 2'd2, 2'd0, 2'd0, 2'd3, 
        2'd2, 2'd1, 2'd1, 2'd0, 2'd2, 2'd3, 2'd2, 2'd2, 
        2'd3, 2'd2, 2'd1, 2'd0, 2'd1, 2'd3, 2'd1, 2'd3, 
        2'd0, 2'd3, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd2, 
        2'd0, 2'd3, 2'd0, 2'd1, 2'd3, 2'd3, 2'd2, 2'd3
        } ),
        .LOC( { 3'd0, 3'd7, 3'd5, 3'd3, 3'd1, 3'd0 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn2_r3_1(
        .din ( din                  ),
        .key ( key[11:6 ]           ),
        .dout( { dout[2], dout[0] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd1, 2'd3, 2'd3, 2'd0, 2'd1, 2'd2, 2'd0, 2'd2, 
        2'd0, 2'd3, 2'd1, 2'd3, 2'd2, 2'd2, 2'd2, 2'd3, 
        2'd1, 2'd2, 2'd3, 2'd2, 2'd0, 2'd3, 2'd1, 2'd0, 
        2'd2, 2'd1, 2'd0, 2'd0, 2'd2, 2'd2, 2'd2, 2'd1, 
        2'd2, 2'd0, 2'd0, 2'd0, 2'd1, 2'd2, 2'd2, 2'd3, 
        2'd3, 2'd0, 2'd3, 2'd0, 2'd3, 2'd1, 2'd3, 2'd2, 
        2'd2, 2'd3, 2'd2, 2'd1, 2'd3, 2'd1, 2'd0, 2'd0, 
        2'd0, 2'd3, 2'd3, 2'd2, 2'd0, 2'd1, 2'd2, 2'd2
        } ),
        .LOC( { 3'd7, 3'd5, 3'd3, 3'd2, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r3_2(
        .din ( din                  ),
        .key ( key[17:12]           ),
        .dout( { dout[6], dout[1] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd1, 2'd1, 2'd2, 2'd2, 2'd0, 2'd3, 2'd2, 2'd0, 
        2'd3, 2'd3, 2'd2, 2'd2, 2'd0, 2'd2, 2'd2, 2'd3, 
        2'd2, 2'd3, 2'd2, 2'd2, 2'd0, 2'd0, 2'd1, 2'd2, 
        2'd1, 2'd1, 2'd1, 2'd2, 2'd0, 2'd1, 2'd3, 2'd3, 
        2'd2, 2'd1, 2'd1, 2'd1, 2'd3, 2'd3, 2'd1, 2'd0, 
        2'd2, 2'd1, 2'd1, 2'd2, 2'd1, 2'd1, 2'd1, 2'd0, 
        2'd0, 2'd2, 2'd2, 2'd1, 2'd1, 2'd0, 2'd1, 2'd3, 
        2'd3, 2'd1, 2'd2, 2'd0, 2'd2, 2'd3, 2'd2, 2'd1
        } ),
        .LOC( { 3'd7, 3'd6, 3'd5, 3'd4, 3'd2, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r3_3(
        .din ( din                  ),
        .key ( key[23:18]           ),
        .dout( { dout[7], dout[4] } )
    );

endmodule


module jtcps2_sbox_fn2_r4(
    input  [ 7:0] din,
    input  [23:0] key,
    output [ 7:0] dout
);

    jtcps2_sbox #(
        .LUT( {
        2'd0, 2'd1, 2'd1, 2'd3, 2'd3, 2'd1, 2'd1, 2'd1, 
        2'd3, 2'd3, 2'd0, 2'd2, 2'd1, 2'd0, 2'd1, 2'd1, 
        2'd1, 2'd3, 2'd2, 2'd1, 2'd1, 2'd0, 2'd0, 2'd2, 
        2'd3, 2'd1, 2'd3, 2'd2, 2'd0, 2'd2, 2'd0, 2'd3, 
        2'd1, 2'd0, 2'd2, 2'd3, 2'd2, 2'd2, 2'd3, 2'd3, 
        2'd2, 2'd0, 2'd3, 2'd2, 2'd0, 2'd2, 2'd1, 2'd0, 
        2'd2, 2'd0, 2'd1, 2'd0, 2'd2, 2'd1, 2'd1, 2'd1, 
        2'd3, 2'd3, 2'd1, 2'd2, 2'd1, 2'd1, 2'd0, 2'd2
        } ),
        .LOC( { 3'd0, 3'd7, 3'd6, 3'd3, 3'd1, 3'd0 } ),
        .OK ( 6'b01_1111 ))
    u_sbox_fn2_r4_0(
        .din ( din                  ),
        .key ( key[ 5:0 ]           ),
        .dout( { dout[3], dout[0] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd2, 2'd0, 2'd1, 2'd2, 2'd3, 2'd1, 2'd2, 2'd3, 
        2'd2, 2'd3, 2'd3, 2'd0, 2'd2, 2'd1, 2'd0, 2'd0, 
        2'd0, 2'd3, 2'd1, 2'd0, 2'd1, 2'd0, 2'd3, 2'd3, 
        2'd3, 2'd1, 2'd3, 2'd2, 2'd2, 2'd1, 2'd2, 2'd2, 
        2'd3, 2'd3, 2'd2, 2'd3, 2'd2, 2'd0, 2'd1, 2'd2, 
        2'd0, 2'd1, 2'd2, 2'd0, 2'd1, 2'd0, 2'd1, 2'd1, 
        2'd0, 2'd1, 2'd0, 2'd1, 2'd2, 2'd2, 2'd2, 2'd0, 
        2'd1, 2'd3, 2'd3, 2'd0, 2'd1, 2'd2, 2'd2, 2'd1
        } ),
        .LOC( { 3'd6, 3'd5, 3'd4, 3'd2, 3'd1, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r4_1(
        .din ( din                  ),
        .key ( key[11:6 ]           ),
        .dout( { dout[7], dout[4] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd3, 2'd1, 2'd1, 2'd2, 2'd3, 2'd0, 2'd0, 2'd1, 
        2'd2, 2'd3, 2'd2, 2'd1, 2'd2, 2'd1, 2'd0, 2'd0, 
        2'd3, 2'd1, 2'd0, 2'd1, 2'd0, 2'd2, 2'd3, 2'd3, 
        2'd1, 2'd1, 2'd3, 2'd0, 2'd0, 2'd1, 2'd3, 2'd0, 
        2'd2, 2'd1, 2'd2, 2'd0, 2'd1, 2'd2, 2'd2, 2'd3, 
        2'd1, 2'd2, 2'd2, 2'd2, 2'd1, 2'd0, 2'd1, 2'd3, 
        2'd2, 2'd3, 2'd0, 2'd0, 2'd1, 2'd1, 2'd2, 2'd0, 
        2'd0, 2'd3, 2'd2, 2'd3, 2'd1, 2'd2, 2'd3, 2'd2
        } ),
        .LOC( { 3'd7, 3'd5, 3'd4, 3'd3, 3'd2, 3'd0 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r4_2(
        .din ( din                  ),
        .key ( key[17:12]           ),
        .dout( { dout[2], dout[1] } )
    );

    jtcps2_sbox #(
        .LUT( {
        2'd1, 2'd2, 2'd3, 2'd1, 2'd0, 2'd0, 2'd3, 2'd2, 
        2'd3, 2'd1, 2'd2, 2'd3, 2'd2, 2'd0, 2'd3, 2'd0, 
        2'd2, 2'd3, 2'd1, 2'd1, 2'd3, 2'd0, 2'd1, 2'd0, 
        2'd3, 2'd3, 2'd1, 2'd2, 2'd2, 2'd0, 2'd3, 2'd1, 
        2'd0, 2'd3, 2'd0, 2'd2, 2'd3, 2'd2, 2'd2, 2'd3, 
        2'd0, 2'd2, 2'd0, 2'd1, 2'd2, 2'd3, 2'd0, 2'd1, 
        2'd3, 2'd0, 2'd0, 2'd2, 2'd1, 2'd1, 2'd3, 2'd3, 
        2'd1, 2'd2, 2'd2, 2'd2, 2'd3, 2'd0, 2'd0, 2'd2
        } ),
        .LOC( { 3'd7, 3'd6, 3'd5, 3'd4, 3'd3, 3'd2 } ),
        .OK ( 6'b11_1111 ))
    u_sbox_fn2_r4_3(
        .din ( din                  ),
        .key ( key[23:18]           ),
        .dout( { dout[6], dout[5] } )
    );

endmodule

