module t48_int
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  [2:0] clk_mstate_i,
   input  jtf_executed_i,
   input  tim_overflow_i,
   input  en_tcnti_i,
   input  dis_tcnti_i,
   input  int_n_i,
   input  ale_i,
   input  last_cycle_i,
   input  en_i_i,
   input  dis_i_i,
   input  retr_executed_i,
   input  int_executed_i,
   output tf_o,
   output ext_int_o,
   output tim_int_o,
   output int_pending_o,
   output int_in_progress_o);
  wire [1:0] int_state_s;
  wire [1:0] int_state_q;
  wire timer_flag_q;
  wire timer_overflow_q;
  wire timer_int_enable_q;
  wire int_q;
  wire int_enable_q;
  wire ale_q;
  wire int_type_q;
  wire int_in_progress_q;
  wire n4944_o;
  wire n4946_o;
  wire n4947_o;
  wire [1:0] n4949_o;
  wire n4951_o;
  wire [1:0] n4953_o;
  wire n4955_o;
  wire [1:0] n4957_o;
  wire n4959_o;
  wire [2:0] n4960_o;
  reg [1:0] n4962_o;
  wire n4965_o;
  wire n4968_o;
  wire n4970_o;
  wire n4971_o;
  wire n4972_o;
  wire n4973_o;
  wire n4974_o;
  wire n4976_o;
  wire n4978_o;
  wire n4980_o;
  wire n4982_o;
  wire n4984_o;
  wire n4986_o;
  wire n4987_o;
  wire n4988_o;
  wire n4989_o;
  wire n4991_o;
  wire n4998_o;
  wire n4999_o;
  wire n5000_o;
  wire n5002_o;
  wire n5003_o;
  wire n5005_o;
  wire n5036_o;
  wire n5038_o;
  wire n5039_o;
  wire n5040_o;
  wire n5048_o;
  wire n5049_o;
  wire n5051_o;
  wire n5067_o;
  wire n5068_o;
  wire n5070_o;
  wire n5072_o;
  wire n5073_o;
  wire [1:0] n5074_o;
  reg [1:0] n5075_q;
  wire n5076_o;
  reg n5077_q;
  wire n5078_o;
  reg n5079_q;
  wire n5080_o;
  reg n5081_q;
  wire n5082_o;
  reg n5083_q;
  wire n5084_o;
  reg n5085_q;
  wire n5086_o;
  reg n5087_q;
  wire n5088_o;
  reg n5089_q;
  wire n5090_o;
  reg n5091_q;
  assign tf_o = n5067_o;
  assign ext_int_o = int_type_q;
  assign tim_int_o = n5068_o;
  assign int_pending_o = n5070_o;
  assign int_in_progress_o = n5073_o;
  /* int.vhd:91:10  */
  assign int_state_s = n4962_o; // (signal)
  /* int.vhd:92:10  */
  assign int_state_q = n5075_q; // (signal)
  /* int.vhd:94:10  */
  assign timer_flag_q = n5077_q; // (signal)
  /* int.vhd:95:10  */
  assign timer_overflow_q = n5079_q; // (signal)
  /* int.vhd:96:10  */
  assign timer_int_enable_q = n5081_q; // (signal)
  /* int.vhd:97:10  */
  assign int_q = n5083_q; // (signal)
  /* int.vhd:98:10  */
  assign int_enable_q = n5085_q; // (signal)
  /* int.vhd:99:10  */
  assign ale_q = n5087_q; // (signal)
  /* int.vhd:100:10  */
  assign int_type_q = n5089_q; // (signal)
  /* int.vhd:101:10  */
  assign int_in_progress_q = n5091_q; // (signal)
  /* int.vhd:123:30  */
  assign n4944_o = last_cycle_i & int_in_progress_q;
  /* int.vhd:124:42  */
  assign n4946_o = clk_mstate_i == 3'b100;
  /* int.vhd:124:25  */
  assign n4947_o = n4946_o & n4944_o;
  /* int.vhd:123:9  */
  assign n4949_o = n4947_o ? 2'b01 : int_state_q;
  /* int.vhd:122:7  */
  assign n4951_o = int_state_q == 2'b00;
  /* int.vhd:129:9  */
  assign n4953_o = int_executed_i ? 2'b10 : int_state_q;
  /* int.vhd:128:7  */
  assign n4955_o = int_state_q == 2'b01;
  /* int.vhd:134:9  */
  assign n4957_o = retr_executed_i ? 2'b00 : int_state_q;
  /* int.vhd:133:7  */
  assign n4959_o = int_state_q == 2'b10;
  assign n4960_o = {n4959_o, n4955_o, n4951_o};
  /* int.vhd:121:5  */
  always @*
    case (n4960_o)
      3'b100: n4962_o = n4957_o;
      3'b010: n4962_o = n4953_o;
      3'b001: n4962_o = n4949_o;
      default: n4962_o = 2'b00;
    endcase
  /* int.vhd:158:14  */
  assign n4965_o = ~res_i;
  /* int.vhd:174:9  */
  assign n4968_o = tim_overflow_i ? 1'b1 : timer_flag_q;
  /* int.vhd:172:9  */
  assign n4970_o = jtf_executed_i ? 1'b0 : n4968_o;
  /* int.vhd:178:24  */
  assign n4971_o = ~int_type_q;
  /* int.vhd:178:36  */
  assign n4972_o = int_executed_i & n4971_o;
  /* int.vhd:179:11  */
  assign n4973_o = ~timer_int_enable_q;
  /* int.vhd:178:56  */
  assign n4974_o = n4972_o | n4973_o;
  /* int.vhd:181:9  */
  assign n4976_o = tim_overflow_i ? 1'b1 : timer_overflow_q;
  /* int.vhd:178:9  */
  assign n4978_o = n4974_o ? 1'b0 : n4976_o;
  /* int.vhd:187:9  */
  assign n4980_o = en_tcnti_i ? 1'b1 : timer_int_enable_q;
  /* int.vhd:185:9  */
  assign n4982_o = dis_tcnti_i ? 1'b0 : n4980_o;
  /* int.vhd:193:9  */
  assign n4984_o = en_i_i ? 1'b1 : int_enable_q;
  /* int.vhd:191:9  */
  assign n4986_o = dis_i_i ? 1'b0 : n4984_o;
  /* int.vhd:199:22  */
  assign n4987_o = int_enable_q & int_q;
  /* int.vhd:199:40  */
  assign n4988_o = n4987_o | timer_overflow_q;
  /* int.vhd:202:14  */
  assign n4989_o = ~int_in_progress_q;
  /* int.vhd:203:45  */
  assign n4991_o = int_enable_q & int_q;
  /* t48_pack-p.vhd:66:5  */
  assign n4998_o = n4991_o ? 1'b1 : 1'b0;
  /* int.vhd:199:9  */
  assign n4999_o = n5000_o ? n4998_o : int_type_q;
  /* int.vhd:199:9  */
  assign n5000_o = n4988_o & n4989_o;
  /* int.vhd:199:9  */
  assign n5002_o = n4988_o ? 1'b1 : int_in_progress_q;
  /* int.vhd:197:9  */
  assign n5003_o = retr_executed_i ? int_type_q : n4999_o;
  /* int.vhd:197:9  */
  assign n5005_o = retr_executed_i ? 1'b0 : n5002_o;
  /* int.vhd:224:14  */
  assign n5036_o = ~res_i;
  /* int.vhd:232:25  */
  assign n5038_o = ale_q & last_cycle_i;
  /* int.vhd:233:22  */
  assign n5039_o = ~ale_i;
  /* int.vhd:233:18  */
  assign n5040_o = n5039_o & n5038_o;
  /* t48_pack-p.vhd:75:5  */
  assign n5048_o = int_n_i ? 1'b1 : 1'b0;
  /* int.vhd:234:20  */
  assign n5049_o = ~n5048_o;
  /* int.vhd:229:7  */
  assign n5051_o = xtal_en_i & n5040_o;
  /* t48_pack-p.vhd:66:5  */
  assign n5067_o = timer_flag_q ? 1'b1 : 1'b0;
  /* int.vhd:249:35  */
  assign n5068_o = ~int_type_q;
  /* int.vhd:250:36  */
  assign n5070_o = int_state_q == 2'b01;
  /* int.vhd:251:58  */
  assign n5072_o = int_state_q != 2'b00;
  /* int.vhd:251:42  */
  assign n5073_o = n5072_o & int_in_progress_q;
  /* int.vhd:167:5  */
  assign n5074_o = en_clk_i ? int_state_s : int_state_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n4965_o)
    if (n4965_o)
      n5075_q <= 2'b00;
    else
      n5075_q <= n5074_o;
  /* int.vhd:167:5  */
  assign n5076_o = en_clk_i ? n4970_o : timer_flag_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n4965_o)
    if (n4965_o)
      n5077_q <= 1'b0;
    else
      n5077_q <= n5076_o;
  /* int.vhd:167:5  */
  assign n5078_o = en_clk_i ? n4978_o : timer_overflow_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n4965_o)
    if (n4965_o)
      n5079_q <= 1'b0;
    else
      n5079_q <= n5078_o;
  /* int.vhd:167:5  */
  assign n5080_o = en_clk_i ? n4982_o : timer_int_enable_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n4965_o)
    if (n4965_o)
      n5081_q <= 1'b0;
    else
      n5081_q <= n5080_o;
  /* int.vhd:228:5  */
  assign n5082_o = n5051_o ? n5049_o : int_q;
  /* int.vhd:228:5  */
  always @(posedge xtal_i or posedge n5036_o)
    if (n5036_o)
      n5083_q <= 1'b0;
    else
      n5083_q <= n5082_o;
  /* int.vhd:167:5  */
  assign n5084_o = en_clk_i ? n4986_o : int_enable_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n4965_o)
    if (n4965_o)
      n5085_q <= 1'b0;
    else
      n5085_q <= n5084_o;
  /* int.vhd:228:5  */
  assign n5086_o = xtal_en_i ? ale_i : ale_q;
  /* int.vhd:228:5  */
  always @(posedge xtal_i or posedge n5036_o)
    if (n5036_o)
      n5087_q <= 1'b0;
    else
      n5087_q <= n5086_o;
  /* int.vhd:167:5  */
  assign n5088_o = en_clk_i ? n5003_o : int_type_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n4965_o)
    if (n4965_o)
      n5089_q <= 1'b0;
    else
      n5089_q <= n5088_o;
  /* int.vhd:167:5  */
  assign n5090_o = en_clk_i ? n5005_o : int_in_progress_q;
  /* int.vhd:167:5  */
  always @(posedge clk_i or posedge n4965_o)
    if (n4965_o)
      n5091_q <= 1'b0;
    else
      n5091_q <= n5090_o;
endmodule

module t48_psw
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  read_psw_i,
   input  read_sp_i,
   input  write_psw_i,
   input  write_sp_i,
   input  special_data_i,
   input  inc_stackp_i,
   input  dec_stackp_i,
   input  write_carry_i,
   input  write_aux_carry_i,
   input  write_f0_i,
   input  write_bs_i,
   input  aux_carry_i,
   output [7:0] data_o,
   output carry_o,
   output aux_carry_o,
   output f0_o,
   output bs_o);
  wire [3:0] psw_q;
  wire [2:0] sp_q;
  wire n4876_o;
  wire [2:0] n4880_o;
  wire [2:0] n4881_o;
  wire [2:0] n4883_o;
  wire [2:0] n4884_o;
  wire [2:0] n4886_o;
  wire [2:0] n4887_o;
  wire n4888_o;
  wire n4889_o;
  wire n4890_o;
  wire n4891_o;
  wire n4895_o;
  wire n4896_o;
  wire n4897_o;
  wire n4898_o;
  wire n4902_o;
  wire n4903_o;
  wire n4904_o;
  wire n4905_o;
  wire n4906_o;
  wire n4907_o;
  wire n4908_o;
  wire n4909_o;
  wire [3:0] n4910_o;
  wire [3:0] n4922_o;
  localparam [7:0] n4923_o = 8'b11111111;
  wire [3:0] n4924_o;
  wire [3:0] n4926_o;
  wire [3:0] n4927_o;
  wire n4929_o;
  wire n4930_o;
  wire n4931_o;
  wire n4932_o;
  wire [3:0] n4933_o;
  reg [3:0] n4934_q;
  wire [2:0] n4935_o;
  reg [2:0] n4936_q;
  wire [7:0] n4937_o;
  assign data_o = n4937_o;
  assign carry_o = n4929_o;
  assign aux_carry_o = n4930_o;
  assign f0_o = n4931_o;
  assign bs_o = n4932_o;
  /* psw.vhd:101:10  */
  assign psw_q = n4934_q; // (signal)
  /* psw.vhd:103:10  */
  assign sp_q = n4936_q; // (signal)
  /* psw.vhd:119:14  */
  assign n4876_o = ~res_i;
  /* psw.vhd:131:34  */
  assign n4880_o = data_i[2:0];
  /* psw.vhd:130:9  */
  assign n4881_o = write_sp_i ? n4880_o : sp_q;
  /* psw.vhd:136:25  */
  assign n4883_o = sp_q + 3'b001;
  /* psw.vhd:135:9  */
  assign n4884_o = inc_stackp_i ? n4883_o : n4881_o;
  /* psw.vhd:140:25  */
  assign n4886_o = sp_q - 3'b001;
  /* psw.vhd:139:9  */
  assign n4887_o = dec_stackp_i ? n4886_o : n4884_o;
  assign n4888_o = data_i[7];
  assign n4889_o = psw_q[3];
  /* psw.vhd:127:9  */
  assign n4890_o = write_psw_i ? n4888_o : n4889_o;
  /* psw.vhd:144:9  */
  assign n4891_o = write_carry_i ? special_data_i : n4890_o;
  assign n4895_o = data_i[6];
  assign n4896_o = psw_q[2];
  /* psw.vhd:127:9  */
  assign n4897_o = write_psw_i ? n4895_o : n4896_o;
  /* psw.vhd:148:9  */
  assign n4898_o = write_aux_carry_i ? aux_carry_i : n4897_o;
  assign n4902_o = data_i[5];
  assign n4903_o = psw_q[1];
  /* psw.vhd:127:9  */
  assign n4904_o = write_psw_i ? n4902_o : n4903_o;
  /* psw.vhd:152:9  */
  assign n4905_o = write_f0_i ? special_data_i : n4904_o;
  assign n4906_o = data_i[4];
  assign n4907_o = psw_q[0];
  /* psw.vhd:127:9  */
  assign n4908_o = write_psw_i ? n4906_o : n4907_o;
  /* psw.vhd:156:9  */
  assign n4909_o = write_bs_i ? special_data_i : n4908_o;
  assign n4910_o = {n4891_o, n4898_o, n4905_o, n4909_o};
  /* psw.vhd:182:5  */
  assign n4922_o = read_psw_i ? psw_q : 4'b1111;
  assign n4924_o = n4923_o[3:0];
  /* psw.vhd:187:33  */
  assign n4926_o = {1'b1, sp_q};
  /* psw.vhd:186:5  */
  assign n4927_o = read_sp_i ? n4926_o : n4924_o;
  /* psw.vhd:207:23  */
  assign n4929_o = psw_q[3];
  /* psw.vhd:208:23  */
  assign n4930_o = psw_q[2];
  /* psw.vhd:209:23  */
  assign n4931_o = psw_q[1];
  /* psw.vhd:210:23  */
  assign n4932_o = psw_q[0];
  /* psw.vhd:123:5  */
  assign n4933_o = en_clk_i ? n4910_o : psw_q;
  /* psw.vhd:123:5  */
  always @(posedge clk_i or posedge n4876_o)
    if (n4876_o)
      n4934_q <= 4'b0000;
    else
      n4934_q <= n4933_o;
  /* psw.vhd:123:5  */
  assign n4935_o = en_clk_i ? n4887_o : sp_q;
  /* psw.vhd:123:5  */
  always @(posedge clk_i or posedge n4876_o)
    if (n4876_o)
      n4936_q <= 3'b000;
    else
      n4936_q <= n4935_o;
  /* psw.vhd:119:5  */
  assign n4937_o = {n4922_o, n4927_o};
endmodule

module t48_pmem_ctrl
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_pcl_i,
   input  read_pcl_i,
   input  write_pch_i,
   input  read_pch_i,
   input  inc_pc_i,
   input  write_pmem_addr_i,
   input  [1:0] addr_type_i,
   input  read_pmem_i,
   input  [7:0] pmem_data_i,
   output [7:0] data_o,
   output [11:0] pmem_addr_o);
  wire [11:0] program_counter_q;
  wire [11:0] pmem_addr_s;
  wire [11:0] pmem_addr_q;
  wire n4802_o;
  wire [3:0] n4804_o;
  wire [10:0] n4805_o;
  wire [10:0] n4807_o;
  wire [10:0] n4808_o;
  wire [10:0] n4809_o;
  wire [7:0] n4810_o;
  wire [7:0] n4811_o;
  wire [7:0] n4812_o;
  wire [2:0] n4813_o;
  wire [2:0] n4814_o;
  wire [2:0] n4815_o;
  wire n4816_o;
  wire n4817_o;
  wire n4818_o;
  wire [11:0] n4819_o;
  wire [7:0] n4820_o;
  wire [7:0] n4821_o;
  wire [3:0] n4822_o;
  wire [3:0] n4823_o;
  wire [3:0] n4824_o;
  wire [11:0] n4826_o;
  wire n4828_o;
  wire n4838_o;
  wire n4840_o;
  wire n4843_o;
  wire [2:0] n4844_o;
  wire [7:0] n4845_o;
  reg [7:0] n4846_o;
  wire [3:0] n4847_o;
  reg [3:0] n4848_o;
  wire [7:0] n4852_o;
  wire [3:0] n4853_o;
  wire [3:0] n4855_o;
  wire [3:0] n4856_o;
  wire [3:0] n4857_o;
  wire [3:0] n4858_o;
  wire [3:0] n4860_o;
  wire [7:0] n4861_o;
  wire [7:0] n4862_o;
  wire [11:0] n4865_o;
  reg [11:0] n4866_q;
  wire [11:0] n4867_o;
  wire [11:0] n4868_o;
  reg [11:0] n4869_q;
  assign data_o = n4862_o;
  assign pmem_addr_o = pmem_addr_q;
  /* pmem_ctrl.vhd:98:10  */
  assign program_counter_q = n4866_q; // (signal)
  /* pmem_ctrl.vhd:102:10  */
  assign pmem_addr_s = n4867_o; // (signal)
  /* pmem_ctrl.vhd:103:10  */
  assign pmem_addr_q = n4869_q; // (signal)
  /* pmem_ctrl.vhd:115:14  */
  assign n4802_o = ~res_i;
  /* pmem_ctrl.vhd:127:28  */
  assign n4804_o = data_i[3:0];
  /* pmem_ctrl.vhd:133:30  */
  assign n4805_o = program_counter_q[10:0];
  /* pmem_ctrl.vhd:133:49  */
  assign n4807_o = n4805_o + 11'b00000000001;
  /* p2.vhd:153:3  */
  assign n4808_o = program_counter_q[10:0];
  /* pmem_ctrl.vhd:128:9  */
  assign n4809_o = inc_pc_i ? n4807_o : n4808_o;
  /* p2.vhd:115:5  */
  assign n4810_o = n4809_o[7:0];
  /* p2.vhd:115:5  */
  assign n4811_o = program_counter_q[7:0];
  /* pmem_ctrl.vhd:125:9  */
  assign n4812_o = write_pch_i ? n4811_o : n4810_o;
  /* decoder.vhd:521:15  */
  assign n4813_o = n4809_o[10:8];
  /* decoder.vhd:521:15  */
  assign n4814_o = n4804_o[2:0];
  /* pmem_ctrl.vhd:125:9  */
  assign n4815_o = write_pch_i ? n4814_o : n4813_o;
  /* p2.vhd:155:5  */
  assign n4816_o = n4804_o[3];
  assign n4817_o = program_counter_q[11];
  /* pmem_ctrl.vhd:125:9  */
  assign n4818_o = write_pch_i ? n4816_o : n4817_o;
  assign n4819_o = {n4818_o, n4815_o, n4812_o};
  /* decoder_pack-p.vhd:115:14  */
  assign n4820_o = n4819_o[7:0];
  /* pmem_ctrl.vhd:123:9  */
  assign n4821_o = write_pcl_i ? data_i : n4820_o;
  /* decoder_pack-p.vhd:114:14  */
  assign n4822_o = n4819_o[11:8];
  assign n4823_o = program_counter_q[11:8];
  /* pmem_ctrl.vhd:123:9  */
  assign n4824_o = write_pcl_i ? n4823_o : n4822_o;
  assign n4826_o = {n4824_o, n4821_o};
  /* pmem_ctrl.vhd:120:7  */
  assign n4828_o = en_clk_i & write_pmem_addr_i;
  /* pmem_ctrl.vhd:165:7  */
  assign n4838_o = addr_type_i == 2'b00;
  /* pmem_ctrl.vhd:169:7  */
  assign n4840_o = addr_type_i == 2'b01;
  /* pmem_ctrl.vhd:175:7  */
  assign n4843_o = addr_type_i == 2'b10;
  assign n4844_o = {n4843_o, n4840_o, n4838_o};
  assign n4845_o = program_counter_q[7:0];
  /* pmem_ctrl.vhd:164:5  */
  always @*
    case (n4844_o)
      3'b100: n4846_o = data_i;
      3'b010: n4846_o = data_i;
      3'b001: n4846_o = n4845_o;
      default: n4846_o = n4845_o;
    endcase
  assign n4847_o = program_counter_q[11:8];
  /* pmem_ctrl.vhd:164:5  */
  always @*
    case (n4844_o)
      3'b100: n4848_o = 4'b0011;
      3'b010: n4848_o = n4847_o;
      3'b001: n4848_o = n4847_o;
      default: n4848_o = n4847_o;
    endcase
  /* pmem_ctrl.vhd:207:51  */
  assign n4852_o = program_counter_q[7:0];
  /* pmem_ctrl.vhd:209:63  */
  assign n4853_o = program_counter_q[11:8];
  /* pmem_ctrl.vhd:208:5  */
  assign n4855_o = read_pch_i ? n4853_o : 4'b1111;
  assign n4856_o = n4852_o[3:0];
  /* pmem_ctrl.vhd:206:5  */
  assign n4857_o = read_pcl_i ? n4856_o : n4855_o;
  assign n4858_o = n4852_o[7:4];
  /* pmem_ctrl.vhd:206:5  */
  assign n4860_o = read_pcl_i ? n4858_o : 4'b1111;
  assign n4861_o = {n4860_o, n4857_o};
  /* pmem_ctrl.vhd:204:5  */
  assign n4862_o = read_pmem_i ? pmem_data_i : n4861_o;
  /* pmem_ctrl.vhd:119:5  */
  assign n4865_o = en_clk_i ? n4826_o : program_counter_q;
  /* pmem_ctrl.vhd:119:5  */
  always @(posedge clk_i or posedge n4802_o)
    if (n4802_o)
      n4866_q <= 12'b000000000000;
    else
      n4866_q <= n4865_o;
  /* pmem_ctrl.vhd:115:5  */
  assign n4867_o = {n4848_o, n4846_o};
  /* pmem_ctrl.vhd:119:5  */
  assign n4868_o = n4828_o ? pmem_addr_s : pmem_addr_q;
  /* pmem_ctrl.vhd:119:5  */
  always @(posedge clk_i or posedge n4802_o)
    if (n4802_o)
      n4869_q <= 12'b000000000000;
    else
      n4869_q <= n4868_o;
endmodule

module t48_p2
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  [7:0] data_i,
   input  write_p2_i,
   input  write_exp_i,
   input  read_p2_i,
   input  read_reg_i,
   input  read_exp_i,
   input  output_pch_i,
   input  [3:0] pch_i,
   input  [7:0] p2_i,
   output [7:0] data_o,
   output [7:0] p2_o,
   output p2l_low_imp_o,
   output p2h_low_imp_o);
  wire [7:0] p2_q;
  wire l_low_imp_q;
  wire h_low_imp_q;
  wire en_clk_q;
  wire l_low_imp_del_q;
  wire h_low_imp_del_q;
  wire output_pch_q;
  wire n4701_o;
  wire [3:0] n4703_o;
  wire [3:0] n4704_o;
  wire [3:0] n4705_o;
  wire n4708_o;
  wire [3:0] n4709_o;
  wire [3:0] n4710_o;
  wire [3:0] n4711_o;
  wire [3:0] n4712_o;
  wire [3:0] n4713_o;
  wire n4715_o;
  wire n4719_o;
  wire [7:0] n4721_o;
  wire n4736_o;
  wire [3:0] n4738_o;
  wire [3:0] n4739_o;
  wire [3:0] n4740_o;
  wire n4741_o;
  wire n4742_o;
  wire n4743_o;
  wire n4746_o;
  wire n4747_o;
  wire n4750_o;
  wire [7:0] n4751_o;
  wire [3:0] n4774_o;
  wire [7:0] n4776_o;
  wire [7:0] n4777_o;
  wire [7:0] n4778_o;
  wire [7:0] n4780_o;
  wire [7:0] n4783_o;
  reg [7:0] n4784_q;
  wire n4785_o;
  reg n4786_q;
  wire n4787_o;
  reg n4788_q;
  wire n4789_o;
  reg n4790_q;
  wire n4791_o;
  reg n4792_q;
  wire n4793_o;
  reg n4794_q;
  wire n4795_o;
  reg n4796_q;
  wire [7:0] n4797_o;
  reg [7:0] n4798_q;
  assign data_o = n4780_o;
  assign p2_o = n4798_q;
  assign p2l_low_imp_o = l_low_imp_del_q;
  assign p2h_low_imp_o = h_low_imp_del_q;
  /* p2.vhd:89:10  */
  assign p2_q = n4784_q; // (signal)
  /* p2.vhd:92:10  */
  assign l_low_imp_q = n4786_q; // (signal)
  /* p2.vhd:93:10  */
  assign h_low_imp_q = n4788_q; // (signal)
  /* p2.vhd:95:10  */
  assign en_clk_q = n4790_q; // (signal)
  /* p2.vhd:96:10  */
  assign l_low_imp_del_q = n4792_q; // (signal)
  /* p2.vhd:97:10  */
  assign h_low_imp_del_q = n4794_q; // (signal)
  /* p2.vhd:98:10  */
  assign output_pch_q = n4796_q; // (signal)
  /* p2.vhd:110:14  */
  assign n4701_o = ~res_i;
  /* p2.vhd:129:41  */
  assign n4703_o = data_i[3:0];
  /* decoder.vhd:496:15  */
  assign n4704_o = p2_q[3:0];
  /* p2.vhd:127:9  */
  assign n4705_o = write_exp_i ? n4703_o : n4704_o;
  /* p2.vhd:127:9  */
  assign n4708_o = write_exp_i ? 1'b1 : 1'b0;
  /* decoder.vhd:521:15  */
  assign n4709_o = data_i[3:0];
  /* p2.vhd:121:9  */
  assign n4710_o = write_p2_i ? n4709_o : n4705_o;
  /* decoder.vhd:521:15  */
  assign n4711_o = data_i[7:4];
  /* decoder.vhd:521:15  */
  assign n4712_o = p2_q[7:4];
  /* p2.vhd:121:9  */
  assign n4713_o = write_p2_i ? n4711_o : n4712_o;
  /* p2.vhd:121:9  */
  assign n4715_o = write_p2_i ? 1'b1 : n4708_o;
  /* p2.vhd:121:9  */
  assign n4719_o = write_p2_i ? 1'b1 : 1'b0;
  assign n4721_o = {n4713_o, n4710_o};
  /* p2.vhd:155:14  */
  assign n4736_o = ~res_i;
  /* decoder.vhd:506:15  */
  assign n4738_o = p2_q[3:0];
  /* p2.vhd:170:9  */
  assign n4739_o = output_pch_i ? pch_i : n4738_o;
  /* decoder.vhd:499:26  */
  assign n4740_o = p2_q[7:4];
  /* p2.vhd:179:26  */
  assign n4741_o = output_pch_q ^ output_pch_i;
  /* p2.vhd:179:44  */
  assign n4742_o = n4741_o | l_low_imp_q;
  /* p2.vhd:178:21  */
  assign n4743_o = n4742_o & en_clk_q;
  /* p2.vhd:178:9  */
  assign n4746_o = n4743_o ? 1'b1 : 1'b0;
  /* p2.vhd:189:21  */
  assign n4747_o = h_low_imp_q & en_clk_q;
  /* p2.vhd:189:9  */
  assign n4750_o = n4747_o ? 1'b1 : 1'b0;
  /* decoder.vhd:499:22  */
  assign n4751_o = {n4740_o, n4739_o};
  /* p2.vhd:221:32  */
  assign n4774_o = p2_i[3:0];
  /* p2.vhd:221:26  */
  assign n4776_o = {4'b0000, n4774_o};
  /* p2.vhd:220:7  */
  assign n4777_o = read_exp_i ? n4776_o : p2_i;
  /* p2.vhd:218:7  */
  assign n4778_o = read_reg_i ? p2_q : n4777_o;
  /* p2.vhd:217:5  */
  assign n4780_o = read_p2_i ? n4778_o : 8'b11111111;
  /* p2.vhd:115:5  */
  assign n4783_o = en_clk_i ? n4721_o : p2_q;
  /* p2.vhd:115:5  */
  always @(posedge clk_i or posedge n4701_o)
    if (n4701_o)
      n4784_q <= 8'b11111111;
    else
      n4784_q <= n4783_o;
  /* p2.vhd:115:5  */
  assign n4785_o = en_clk_i ? n4715_o : l_low_imp_q;
  /* p2.vhd:115:5  */
  always @(posedge clk_i or posedge n4701_o)
    if (n4701_o)
      n4786_q <= 1'b0;
    else
      n4786_q <= n4785_o;
  /* p2.vhd:115:5  */
  assign n4787_o = en_clk_i ? n4719_o : h_low_imp_q;
  /* p2.vhd:115:5  */
  always @(posedge clk_i or posedge n4701_o)
    if (n4701_o)
      n4788_q <= 1'b0;
    else
      n4788_q <= n4787_o;
  /* p2.vhd:162:5  */
  assign n4789_o = xtal_en_i ? en_clk_i : en_clk_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4736_o)
    if (n4736_o)
      n4790_q <= 1'b0;
    else
      n4790_q <= n4789_o;
  /* p2.vhd:162:5  */
  assign n4791_o = xtal_en_i ? n4746_o : l_low_imp_del_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4736_o)
    if (n4736_o)
      n4792_q <= 1'b0;
    else
      n4792_q <= n4791_o;
  /* p2.vhd:162:5  */
  assign n4793_o = xtal_en_i ? n4750_o : h_low_imp_del_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4736_o)
    if (n4736_o)
      n4794_q <= 1'b0;
    else
      n4794_q <= n4793_o;
  /* p2.vhd:162:5  */
  assign n4795_o = xtal_en_i ? output_pch_i : output_pch_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4736_o)
    if (n4736_o)
      n4796_q <= 1'b0;
    else
      n4796_q <= n4795_o;
  /* p2.vhd:162:5  */
  assign n4797_o = xtal_en_i ? n4751_o : n4798_q;
  /* p2.vhd:162:5  */
  always @(posedge xtal_i or posedge n4736_o)
    if (n4736_o)
      n4798_q <= 8'b11111111;
    else
      n4798_q <= n4797_o;
endmodule

module t48_p1
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_p1_i,
   input  read_p1_i,
   input  read_reg_i,
   input  [7:0] p1_i,
   output [7:0] data_o,
   output [7:0] p1_o,
   output p1_low_imp_o);
  wire [7:0] p1_q;
  wire low_imp_q;
  wire n4671_o;
  wire n4676_o;
  wire n4677_o;
  wire [7:0] n4687_o;
  wire [7:0] n4689_o;
  wire [7:0] n4692_o;
  reg [7:0] n4693_q;
  wire n4694_o;
  reg n4695_q;
  assign data_o = n4689_o;
  assign p1_o = p1_q;
  assign p1_low_imp_o = low_imp_q;
  /* p1.vhd:81:10  */
  assign p1_q = n4693_q; // (signal)
  /* p1.vhd:84:10  */
  assign low_imp_q = n4695_q; // (signal)
  /* p1.vhd:96:14  */
  assign n4671_o = ~res_i;
  /* p1.vhd:103:9  */
  assign n4676_o = write_p1_i ? 1'b1 : 1'b0;
  /* p1.vhd:101:7  */
  assign n4677_o = en_clk_i & write_p1_i;
  /* p1.vhd:133:7  */
  assign n4687_o = read_reg_i ? p1_q : p1_i;
  /* p1.vhd:132:5  */
  assign n4689_o = read_p1_i ? n4687_o : 8'b11111111;
  /* p1.vhd:100:5  */
  assign n4692_o = n4677_o ? data_i : p1_q;
  /* p1.vhd:100:5  */
  always @(posedge clk_i or posedge n4671_o)
    if (n4671_o)
      n4693_q <= 8'b11111111;
    else
      n4693_q <= n4692_o;
  /* p1.vhd:100:5  */
  assign n4694_o = en_clk_i ? n4676_o : low_imp_q;
  /* p1.vhd:100:5  */
  always @(posedge clk_i or posedge n4671_o)
    if (n4671_o)
      n4695_q <= 1'b0;
    else
      n4695_q <= n4694_o;
endmodule

module t48_timer_4
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  t1_i,
   input  [2:0] clk_mstate_i,
   input  [7:0] data_i,
   input  read_timer_i,
   input  write_timer_i,
   input  start_t_i,
   input  start_cnt_i,
   input  stop_tcnt_i,
   output [7:0] data_o,
   output overflow_o);
  wire [7:0] counter_q;
  wire overflow_q;
  wire increment_s;
  wire [1:0] inc_sel_q;
  wire t1_q;
  wire t1_inc_s;
  wire [4:0] prescaler_q;
  wire pre_inc_s;
  wire n4557_o;
  wire n4559_o;
  wire n4561_o;
  wire n4562_o;
  wire n4563_o;
  wire n4566_o;
  wire n4568_o;
  wire n4572_o;
  wire n4574_o;
  wire n4575_o;
  wire n4578_o;
  wire n4580_o;
  wire n4582_o;
  wire [2:0] n4583_o;
  reg n4586_o;
  wire n4590_o;
  wire [7:0] n4593_o;
  wire n4595_o;
  wire n4598_o;
  wire [7:0] n4599_o;
  wire n4601_o;
  wire [7:0] n4602_o;
  wire n4604_o;
  wire n4607_o;
  wire n4609_o;
  wire n4611_o;
  wire n4614_o;
  wire [4:0] n4616_o;
  wire [4:0] n4617_o;
  wire [4:0] n4619_o;
  wire [1:0] n4621_o;
  wire [1:0] n4623_o;
  wire [1:0] n4625_o;
  wire n4629_o;
  wire [7:0] n4647_o;
  wire n4656_o;
  wire [7:0] n4657_o;
  reg [7:0] n4658_q;
  wire n4659_o;
  reg n4660_q;
  wire [1:0] n4661_o;
  reg [1:0] n4662_q;
  wire n4663_o;
  reg n4664_q;
  wire [4:0] n4665_o;
  reg [4:0] n4666_q;
  assign data_o = n4647_o;
  assign overflow_o = n4656_o;
  /* timer.vhd:89:10  */
  assign counter_q = n4658_q; // (signal)
  /* timer.vhd:90:10  */
  assign overflow_q = n4660_q; // (signal)
  /* timer.vhd:94:10  */
  assign increment_s = n4586_o; // (signal)
  /* timer.vhd:95:10  */
  assign inc_sel_q = n4662_q; // (signal)
  /* timer.vhd:98:10  */
  assign t1_q = n4664_q; // (signal)
  /* timer.vhd:99:10  */
  assign t1_inc_s = n4568_o; // (signal)
  /* timer.vhd:102:10  */
  assign prescaler_q = n4666_q; // (signal)
  /* timer.vhd:103:10  */
  assign pre_inc_s = n4575_o; // (signal)
  /* timer.vhd:134:48  */
  assign n4557_o = clk_mstate_i == 3'b011;
  /* timer.vhd:134:31  */
  assign n4559_o = n4557_o & 1'b1;
  /* timer.vhd:133:59  */
  assign n4561_o = 1'b0 | n4559_o;
  /* timer.vhd:136:30  */
  assign n4562_o = ~t1_i;
  /* timer.vhd:136:21  */
  assign n4563_o = n4562_o & t1_q;
  /* timer.vhd:136:7  */
  assign n4566_o = n4563_o ? 1'b1 : 1'b0;
  /* timer.vhd:133:5  */
  assign n4568_o = n4561_o ? n4566_o : 1'b0;
  /* timer.vhd:146:29  */
  assign n4572_o = clk_mstate_i == 3'b011;
  /* timer.vhd:146:55  */
  assign n4574_o = prescaler_q == 5'b11111;
  /* timer.vhd:146:39  */
  assign n4575_o = n4574_o & n4572_o;
  /* timer.vhd:163:7  */
  assign n4578_o = inc_sel_q == 2'b00;
  /* timer.vhd:165:7  */
  assign n4580_o = inc_sel_q == 2'b01;
  /* timer.vhd:167:7  */
  assign n4582_o = inc_sel_q == 2'b10;
  assign n4583_o = {n4582_o, n4580_o, n4578_o};
  /* timer.vhd:162:5  */
  always @*
    case (n4583_o)
      3'b100: n4586_o = t1_inc_s;
      3'b010: n4586_o = pre_inc_s;
      3'b001: n4586_o = 1'b0;
      default: n4586_o = 1'b0;
    endcase
  /* timer.vhd:186:14  */
  assign n4590_o = ~res_i;
  /* timer.vhd:203:37  */
  assign n4593_o = counter_q + 8'b00000001;
  /* timer.vhd:205:24  */
  assign n4595_o = counter_q == 8'b11111111;
  /* timer.vhd:205:11  */
  assign n4598_o = n4595_o ? 1'b1 : 1'b0;
  /* timer.vhd:202:9  */
  assign n4599_o = increment_s ? n4593_o : counter_q;
  /* timer.vhd:202:9  */
  assign n4601_o = increment_s ? n4598_o : 1'b0;
  /* timer.vhd:199:9  */
  assign n4602_o = write_timer_i ? data_i : n4599_o;
  /* timer.vhd:199:9  */
  assign n4604_o = write_timer_i ? 1'b0 : n4601_o;
  /* timer.vhd:213:52  */
  assign n4607_o = clk_mstate_i == 3'b011;
  /* timer.vhd:213:35  */
  assign n4609_o = n4607_o & 1'b1;
  /* timer.vhd:212:63  */
  assign n4611_o = 1'b0 | n4609_o;
  /* timer.vhd:221:28  */
  assign n4614_o = clk_mstate_i == 3'b010;
  /* timer.vhd:222:39  */
  assign n4616_o = prescaler_q + 5'b00001;
  /* timer.vhd:221:9  */
  assign n4617_o = n4614_o ? n4616_o : prescaler_q;
  /* timer.vhd:218:9  */
  assign n4619_o = start_t_i ? 5'b00000 : n4617_o;
  /* timer.vhd:231:9  */
  assign n4621_o = stop_tcnt_i ? 2'b00 : inc_sel_q;
  /* timer.vhd:229:9  */
  assign n4623_o = start_cnt_i ? 2'b10 : n4621_o;
  /* timer.vhd:227:9  */
  assign n4625_o = start_t_i ? 2'b01 : n4623_o;
  /* timer.vhd:194:7  */
  assign n4629_o = en_clk_i & n4611_o;
  /* timer.vhd:248:17  */
  assign n4647_o = read_timer_i ? counter_q : 8'b11111111;
  /* t48_pack-p.vhd:66:5  */
  assign n4656_o = overflow_q ? 1'b1 : 1'b0;
  /* timer.vhd:193:5  */
  assign n4657_o = en_clk_i ? n4602_o : counter_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4590_o)
    if (n4590_o)
      n4658_q <= 8'b00000000;
    else
      n4658_q <= n4657_o;
  /* timer.vhd:193:5  */
  assign n4659_o = en_clk_i ? n4604_o : overflow_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4590_o)
    if (n4590_o)
      n4660_q <= 1'b0;
    else
      n4660_q <= n4659_o;
  /* timer.vhd:193:5  */
  assign n4661_o = en_clk_i ? n4625_o : inc_sel_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4590_o)
    if (n4590_o)
      n4662_q <= 2'b00;
    else
      n4662_q <= n4661_o;
  /* timer.vhd:193:5  */
  assign n4663_o = n4629_o ? t1_i : t1_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4590_o)
    if (n4590_o)
      n4664_q <= 1'b0;
    else
      n4664_q <= n4663_o;
  /* timer.vhd:193:5  */
  assign n4665_o = en_clk_i ? n4619_o : prescaler_q;
  /* timer.vhd:193:5  */
  always @(posedge clk_i or posedge n4590_o)
    if (n4590_o)
      n4666_q <= 5'b00000;
    else
      n4666_q <= n4665_o;
endmodule

module t48_dmem_ctrl
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_dmem_addr_i,
   input  write_dmem_i,
   input  read_dmem_i,
   input  [1:0] addr_type_i,
   input  bank_select_i,
   input  [7:0] dmem_data_i,
   output [7:0] data_o,
   output [7:0] dmem_addr_o,
   output dmem_we_o,
   output [7:0] dmem_data_o);
  wire [7:0] dmem_addr_s;
  wire [7:0] dmem_addr_q;
  wire n4474_o;
  wire [2:0] n4475_o;
  localparam [7:0] n4476_o = 8'b00000000;
  wire [1:0] n4479_o;
  wire [1:0] n4480_o;
  wire [2:0] n4481_o;
  wire n4483_o;
  wire [2:0] n4484_o;
  wire [5:0] n4487_o;
  wire [5:0] n4489_o;
  localparam [7:0] n4490_o = 8'b00000000;
  wire [1:0] n4491_o;
  wire n4493_o;
  wire n4496_o;
  wire [3:0] n4497_o;
  wire n4498_o;
  wire n4499_o;
  wire n4500_o;
  wire n4501_o;
  reg n4502_o;
  wire [1:0] n4503_o;
  wire [1:0] n4504_o;
  wire [1:0] n4505_o;
  wire [1:0] n4506_o;
  reg [1:0] n4507_o;
  wire [1:0] n4508_o;
  wire [1:0] n4509_o;
  wire [1:0] n4510_o;
  reg [1:0] n4511_o;
  wire n4512_o;
  wire n4513_o;
  wire n4514_o;
  wire n4515_o;
  reg n4516_o;
  wire [1:0] n4517_o;
  wire [1:0] n4518_o;
  wire [1:0] n4519_o;
  reg [1:0] n4520_o;
  wire n4530_o;
  wire n4533_o;
  wire n4538_o;
  wire [7:0] n4539_o;
  wire [7:0] n4540_o;
  wire n4549_o;
  wire [7:0] n4550_o;
  wire [7:0] n4551_o;
  reg [7:0] n4552_q;
  assign data_o = n4540_o;
  assign dmem_addr_o = n4539_o;
  assign dmem_we_o = n4549_o;
  assign dmem_data_o = data_i;
  /* dmem_ctrl.vhd:91:10  */
  assign dmem_addr_s = n4550_o; // (signal)
  /* dmem_ctrl.vhd:92:10  */
  assign dmem_addr_q = n4552_q; // (signal)
  /* dmem_ctrl.vhd:112:7  */
  assign n4474_o = addr_type_i == 2'b00;
  /* dmem_ctrl.vhd:117:44  */
  assign n4475_o = data_i[2:0];
  /* decoder.vhd:155:5  */
  assign n4479_o = n4476_o[4:3];
  /* dmem_ctrl.vhd:119:9  */
  assign n4480_o = bank_select_i ? 2'b11 : n4479_o;
  /* decoder.vhd:153:5  */
  assign n4481_o = n4476_o[7:5];
  /* dmem_ctrl.vhd:115:7  */
  assign n4483_o = addr_type_i == 2'b01;
  /* dmem_ctrl.vhd:126:53  */
  assign n4484_o = data_i[2:0];
  /* decoder.vhd:142:5  */
  assign n4487_o = {2'b00, n4484_o, 1'b0};
  /* dmem_ctrl.vhd:128:51  */
  assign n4489_o = n4487_o + 6'b001000;
  /* decoder.vhd:135:5  */
  assign n4491_o = n4490_o[7:6];
  /* dmem_ctrl.vhd:124:7  */
  assign n4493_o = addr_type_i == 2'b10;
  /* dmem_ctrl.vhd:133:7  */
  assign n4496_o = addr_type_i == 2'b11;
  /* decoder.vhd:125:5  */
  assign n4497_o = {n4496_o, n4493_o, n4483_o, n4474_o};
  /* decoder.vhd:124:5  */
  assign n4498_o = data_i[0];
  /* decoder.vhd:123:5  */
  assign n4499_o = n4475_o[0];
  /* decoder.vhd:121:5  */
  assign n4500_o = n4489_o[0];
  /* decoder.vhd:120:5  */
  assign n4501_o = dmem_addr_q[0];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4497_o)
      4'b1000: n4502_o = 1'b1;
      4'b0100: n4502_o = n4500_o;
      4'b0010: n4502_o = n4499_o;
      4'b0001: n4502_o = n4498_o;
      default: n4502_o = n4501_o;
    endcase
  /* decoder.vhd:116:5  */
  assign n4503_o = data_i[2:1];
  /* decoder.vhd:115:5  */
  assign n4504_o = n4475_o[2:1];
  /* decoder.vhd:114:5  */
  assign n4505_o = n4489_o[2:1];
  /* decoder.vhd:113:5  */
  assign n4506_o = dmem_addr_q[2:1];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4497_o)
      4'b1000: n4507_o = n4506_o;
      4'b0100: n4507_o = n4505_o;
      4'b0010: n4507_o = n4504_o;
      4'b0001: n4507_o = n4503_o;
      default: n4507_o = n4506_o;
    endcase
  /* decoder.vhd:109:5  */
  assign n4508_o = data_i[4:3];
  /* decoder.vhd:108:5  */
  assign n4509_o = n4489_o[4:3];
  /* decoder.vhd:107:5  */
  assign n4510_o = dmem_addr_q[4:3];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4497_o)
      4'b1000: n4511_o = n4510_o;
      4'b0100: n4511_o = n4509_o;
      4'b0010: n4511_o = n4480_o;
      4'b0001: n4511_o = n4508_o;
      default: n4511_o = n4510_o;
    endcase
  /* decoder.vhd:105:5  */
  assign n4512_o = data_i[5];
  /* decoder.vhd:104:5  */
  assign n4513_o = n4481_o[0];
  /* decoder.vhd:103:5  */
  assign n4514_o = n4489_o[5];
  /* decoder.vhd:102:5  */
  assign n4515_o = dmem_addr_q[5];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4497_o)
      4'b1000: n4516_o = n4515_o;
      4'b0100: n4516_o = n4514_o;
      4'b0010: n4516_o = n4513_o;
      4'b0001: n4516_o = n4512_o;
      default: n4516_o = n4515_o;
    endcase
  /* decoder.vhd:100:5  */
  assign n4517_o = data_i[7:6];
  /* decoder.vhd:99:5  */
  assign n4518_o = n4481_o[2:1];
  /* decoder.vhd:98:5  */
  assign n4519_o = dmem_addr_q[7:6];
  /* dmem_ctrl.vhd:111:5  */
  always @*
    case (n4497_o)
      4'b1000: n4520_o = n4519_o;
      4'b0100: n4520_o = n4491_o;
      4'b0010: n4520_o = n4518_o;
      4'b0001: n4520_o = n4517_o;
      default: n4520_o = n4519_o;
    endcase
  /* dmem_ctrl.vhd:165:14  */
  assign n4530_o = ~res_i;
  /* dmem_ctrl.vhd:169:7  */
  assign n4533_o = en_clk_i & write_dmem_addr_i;
  /* dmem_ctrl.vhd:188:41  */
  assign n4538_o = en_clk_i & write_dmem_addr_i;
  /* dmem_ctrl.vhd:188:18  */
  assign n4539_o = n4538_o ? dmem_addr_s : dmem_addr_q;
  /* dmem_ctrl.vhd:196:18  */
  assign n4540_o = read_dmem_i ? dmem_data_i : 8'b11111111;
  /* t48_pack-p.vhd:66:5  */
  assign n4549_o = write_dmem_i ? 1'b1 : 1'b0;
  assign n4550_o = {n4520_o, n4516_o, n4511_o, n4507_o, n4502_o};
  /* dmem_ctrl.vhd:168:5  */
  assign n4551_o = n4533_o ? dmem_addr_s : dmem_addr_q;
  /* dmem_ctrl.vhd:168:5  */
  always @(posedge clk_i or posedge n4530_o)
    if (n4530_o)
      n4552_q <= 8'b00000000;
    else
      n4552_q <= n4551_o;
endmodule

module t48_decoder_1_0_0
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  ea_i,
   input  ale_i,
   input  int_n_i,
   input  [7:0] data_i,
   input  bus_set_f1_i,
   input  bus_clear_f1_i,
   input  alu_carry_i,
   input  alu_da_overflow_i,
   input  [2:0] clk_mstate_i,
   input  clk_second_cycle_i,
   input  cnd_take_branch_i,
   input  psw_carry_i,
   input  psw_aux_carry_i,
   input  psw_f0_i,
   input  tim_overflow_i,
   output t0_dir_o,
   output [7:0] data_o,
   output alu_write_accu_o,
   output alu_write_shadow_o,
   output alu_write_temp_reg_o,
   output alu_read_alu_o,
   output bus_write_bus_o,
   output bus_read_bus_o,
   output bus_ibf_int_o,
   output bus_en_dma_o,
   output bus_en_flags_o,
   output bus_write_sts_o,
   output dm_write_dmem_addr_o,
   output dm_write_dmem_o,
   output dm_read_dmem_o,
   output p1_write_p1_o,
   output p1_read_p1_o,
   output p2_write_p2_o,
   output p2_write_exp_o,
   output p2_read_p2_o,
   output p2_read_exp_o,
   output pm_write_pcl_o,
   output pm_read_pcl_o,
   output pm_write_pch_o,
   output pm_read_pch_o,
   output pm_read_pmem_o,
   output psw_read_psw_o,
   output psw_read_sp_o,
   output psw_write_psw_o,
   output psw_write_sp_o,
   output [3:0] alu_op_o,
   output alu_use_carry_o,
   output alu_da_high_o,
   output alu_accu_low_o,
   output alu_p06_temp_reg_o,
   output alu_p60_temp_reg_o,
   output bus_output_pcl_o,
   output bus_bidir_bus_o,
   output clk_multi_cycle_o,
   output clk_assert_psen_o,
   output clk_assert_prog_o,
   output clk_assert_rd_o,
   output clk_assert_wr_o,
   output cnd_compute_take_o,
   output [3:0] cnd_branch_cond_o,
   output [2:0] cnd_comp_value_o,
   output cnd_f1_o,
   output cnd_tf_o,
   output [1:0] dm_addr_type_o,
   output p1_read_reg_o,
   output p2_read_reg_o,
   output p2_output_pch_o,
   output pm_inc_pc_o,
   output pm_write_pmem_addr_o,
   output [1:0] pm_addr_type_o,
   output psw_special_data_o,
   output psw_inc_stackp_o,
   output psw_dec_stackp_o,
   output psw_write_carry_o,
   output psw_write_aux_carry_o,
   output psw_write_f0_o,
   output psw_write_bs_o,
   output tim_read_timer_o,
   output tim_write_timer_o,
   output tim_start_t_o,
   output tim_start_cnt_o,
   output tim_stop_tcnt_o);
  wire opc_multi_cycle_s;
  wire opc_read_bus_s;
  wire opc_inj_int_s;
  wire [7:0] opc_opcode_q;
  wire [5:0] opc_mnemonic_s;
  wire last_cycle_s;
  wire assert_psen_s;
  wire branch_taken_s;
  wire branch_taken_q;
  wire pm_inc_pc_s;
  wire pm_write_pmem_addr_s;
  wire add_inc_pc_s;
  wire add_write_pmem_addr_s;
  wire clear_f1_s;
  wire cpl_f1_s;
  wire f1_q;
  wire clear_mb_s;
  wire set_mb_s;
  wire mb_q;
  wire ent0_clk_s;
  wire t0_dir_q;
  wire [7:0] data_s;
  wire read_dec_s;
  wire tf_s;
  wire bus_read_bus_s;
  wire add_read_bus_s;
  wire dm_write_dmem_s;
  wire p2_output_exp_s;
  wire movx_first_cycle_s;
  wire jtf_executed_s;
  wire en_tcnti_s;
  wire dis_tcnti_s;
  wire en_i_s;
  wire dis_i_s;
  wire tim_int_s;
  wire retr_executed_s;
  wire int_executed_s;
  wire int_pending_s;
  wire int_in_progress_s;
  wire [6:0] mnemonic_rec_s;
  wire [5:0] mnemonic_q;
  wire n1116_o;
  wire n1118_o;
  wire n1119_o;
  wire n1121_o;
  wire n1122_o;
  wire n1124_o;
  wire n1126_o;
  wire n1128_o;
  wire n1130_o;
  wire n1132_o;
  wire n1133_o;
  wire n1135_o;
  wire n1136_o;
  wire n1138_o;
  wire n1139_o;
  wire n1141_o;
  wire n1143_o;
  wire n1144_o;
  wire n1146_o;
  wire n1147_o;
  wire n1149_o;
  wire n1151_o;
  wire n1152_o;
  wire n1154_o;
  wire n1155_o;
  wire n1157_o;
  wire n1159_o;
  wire n1160_o;
  wire [7:0] n1161_o;
  reg [5:0] n1171_o;
  reg n1180_o;
  wire n1183_o;
  wire n1193_o;
  wire n1195_o;
  wire n1196_o;
  wire n1198_o;
  wire n1199_o;
  wire n1201_o;
  wire n1202_o;
  wire n1204_o;
  wire n1205_o;
  wire n1207_o;
  wire n1208_o;
  wire n1210_o;
  wire n1211_o;
  wire n1213_o;
  wire n1214_o;
  wire n1216_o;
  wire n1217_o;
  wire n1219_o;
  wire n1220_o;
  wire n1222_o;
  wire n1223_o;
  wire n1225_o;
  wire n1226_o;
  wire n1228_o;
  wire n1229_o;
  wire n1231_o;
  wire n1232_o;
  wire n1234_o;
  wire n1235_o;
  wire n1237_o;
  wire n1238_o;
  wire n1240_o;
  wire n1241_o;
  wire n1243_o;
  wire n1244_o;
  wire n1246_o;
  wire n1247_o;
  wire n1249_o;
  wire n1250_o;
  wire n1252_o;
  wire n1254_o;
  wire n1255_o;
  wire n1257_o;
  wire n1259_o;
  wire n1260_o;
  wire n1262_o;
  wire n1263_o;
  wire n1265_o;
  wire n1266_o;
  wire n1268_o;
  wire n1269_o;
  wire n1271_o;
  wire n1272_o;
  wire n1274_o;
  wire n1275_o;
  wire n1277_o;
  wire n1278_o;
  wire n1280_o;
  wire n1281_o;
  wire n1283_o;
  wire n1284_o;
  wire n1286_o;
  wire n1288_o;
  wire n1290_o;
  wire n1291_o;
  wire n1293_o;
  wire n1294_o;
  wire n1296_o;
  wire n1297_o;
  wire n1299_o;
  wire n1300_o;
  wire n1302_o;
  wire n1303_o;
  wire n1305_o;
  wire n1306_o;
  wire n1308_o;
  wire n1309_o;
  wire n1311_o;
  wire n1313_o;
  wire n1315_o;
  wire n1317_o;
  wire n1318_o;
  wire n1320_o;
  wire n1322_o;
  wire n1324_o;
  wire n1326_o;
  wire n1327_o;
  wire n1329_o;
  wire n1331_o;
  wire n1333_o;
  wire n1334_o;
  wire n1336_o;
  wire n1337_o;
  wire n1339_o;
  wire n1340_o;
  wire n1342_o;
  wire n1343_o;
  wire n1345_o;
  wire n1346_o;
  wire n1348_o;
  wire n1349_o;
  wire n1351_o;
  wire n1352_o;
  wire n1354_o;
  wire n1355_o;
  wire n1357_o;
  wire n1359_o;
  wire n1360_o;
  wire n1362_o;
  wire n1364_o;
  wire n1365_o;
  wire n1367_o;
  wire n1369_o;
  wire n1370_o;
  wire n1372_o;
  wire n1373_o;
  wire n1375_o;
  wire n1376_o;
  wire n1378_o;
  wire n1379_o;
  wire n1381_o;
  wire n1382_o;
  wire n1384_o;
  wire n1385_o;
  wire n1387_o;
  wire n1388_o;
  wire n1390_o;
  wire n1392_o;
  wire n1393_o;
  wire n1395_o;
  wire n1397_o;
  wire n1398_o;
  wire n1400_o;
  wire n1401_o;
  wire n1403_o;
  wire n1404_o;
  wire n1406_o;
  wire n1407_o;
  wire n1409_o;
  wire n1410_o;
  wire n1412_o;
  wire n1413_o;
  wire n1415_o;
  wire n1416_o;
  wire n1418_o;
  wire n1419_o;
  wire n1421_o;
  wire n1422_o;
  wire n1424_o;
  wire n1425_o;
  wire n1427_o;
  wire n1429_o;
  wire n1430_o;
  wire n1432_o;
  wire n1433_o;
  wire n1435_o;
  wire n1436_o;
  wire n1438_o;
  wire n1439_o;
  wire n1441_o;
  wire n1442_o;
  wire n1444_o;
  wire n1445_o;
  wire n1447_o;
  wire n1448_o;
  wire n1450_o;
  wire n1452_o;
  wire n1453_o;
  wire n1455_o;
  wire n1457_o;
  wire n1458_o;
  wire n1460_o;
  wire n1462_o;
  wire n1463_o;
  wire n1465_o;
  wire n1466_o;
  wire n1468_o;
  wire n1469_o;
  wire n1471_o;
  wire n1472_o;
  wire n1474_o;
  wire n1475_o;
  wire n1477_o;
  wire n1478_o;
  wire n1480_o;
  wire n1481_o;
  wire n1483_o;
  wire n1485_o;
  wire n1487_o;
  wire n1488_o;
  wire n1490_o;
  wire n1491_o;
  wire n1493_o;
  wire n1494_o;
  wire n1496_o;
  wire n1498_o;
  wire n1500_o;
  wire n1501_o;
  wire n1503_o;
  wire n1505_o;
  wire n1507_o;
  wire n1509_o;
  wire n1510_o;
  wire n1512_o;
  wire n1513_o;
  wire n1515_o;
  wire n1516_o;
  wire n1518_o;
  wire n1519_o;
  wire n1521_o;
  wire n1522_o;
  wire n1524_o;
  wire n1525_o;
  wire n1527_o;
  wire n1528_o;
  wire n1530_o;
  wire n1531_o;
  wire n1533_o;
  wire n1534_o;
  wire n1536_o;
  wire n1538_o;
  wire n1540_o;
  wire n1541_o;
  wire n1543_o;
  wire n1544_o;
  wire n1546_o;
  wire n1547_o;
  wire n1549_o;
  wire n1550_o;
  wire n1552_o;
  wire n1553_o;
  wire n1555_o;
  wire n1556_o;
  wire n1558_o;
  wire n1559_o;
  wire n1561_o;
  wire n1562_o;
  wire n1564_o;
  wire n1565_o;
  wire n1567_o;
  wire n1569_o;
  wire n1570_o;
  wire n1572_o;
  wire n1573_o;
  wire n1575_o;
  wire n1576_o;
  wire n1578_o;
  wire n1579_o;
  wire n1581_o;
  wire n1582_o;
  wire n1584_o;
  wire n1585_o;
  wire n1587_o;
  wire n1588_o;
  wire n1590_o;
  wire n1591_o;
  wire n1593_o;
  wire n1594_o;
  wire n1596_o;
  wire n1598_o;
  wire n1599_o;
  wire n1601_o;
  wire n1603_o;
  wire n1604_o;
  wire n1606_o;
  wire n1607_o;
  wire n1609_o;
  wire n1610_o;
  wire n1612_o;
  wire n1614_o;
  wire n1615_o;
  wire n1617_o;
  wire n1619_o;
  wire n1621_o;
  wire n1622_o;
  wire n1624_o;
  wire n1625_o;
  wire n1627_o;
  wire n1628_o;
  wire n1630_o;
  wire n1631_o;
  wire n1633_o;
  wire n1634_o;
  wire n1636_o;
  wire n1637_o;
  wire n1639_o;
  wire n1640_o;
  wire n1642_o;
  wire n1643_o;
  wire n1645_o;
  wire n1646_o;
  wire n1648_o;
  wire n1650_o;
  wire n1652_o;
  wire n1653_o;
  wire n1655_o;
  wire n1656_o;
  wire n1658_o;
  wire n1659_o;
  wire n1661_o;
  wire n1662_o;
  wire n1664_o;
  wire n1665_o;
  wire n1667_o;
  wire n1668_o;
  wire n1670_o;
  wire n1671_o;
  wire n1673_o;
  wire n1674_o;
  wire n1676_o;
  wire n1677_o;
  wire n1679_o;
  wire n1680_o;
  wire n1682_o;
  wire n1683_o;
  wire n1685_o;
  wire n1687_o;
  wire n1688_o;
  wire n1690_o;
  wire n1692_o;
  wire n1693_o;
  wire n1695_o;
  wire n1697_o;
  wire n1698_o;
  wire n1700_o;
  wire n1702_o;
  wire n1703_o;
  wire n1705_o;
  wire n1707_o;
  wire n1709_o;
  wire n1710_o;
  wire n1712_o;
  wire n1714_o;
  wire n1716_o;
  wire n1717_o;
  wire n1719_o;
  wire n1720_o;
  wire n1722_o;
  wire n1723_o;
  wire n1725_o;
  wire n1726_o;
  wire n1728_o;
  wire n1729_o;
  wire n1731_o;
  wire n1732_o;
  wire n1734_o;
  wire n1735_o;
  wire n1737_o;
  wire n1738_o;
  wire n1740_o;
  wire n1741_o;
  wire n1743_o;
  wire n1744_o;
  wire n1746_o;
  wire n1747_o;
  wire n1749_o;
  wire n1751_o;
  wire n1752_o;
  wire n1754_o;
  wire n1755_o;
  wire n1757_o;
  wire n1758_o;
  wire n1760_o;
  wire n1761_o;
  wire n1763_o;
  wire n1764_o;
  wire n1766_o;
  wire n1767_o;
  wire n1769_o;
  wire n1770_o;
  wire n1772_o;
  wire n1773_o;
  wire n1775_o;
  wire n1776_o;
  wire n1778_o;
  wire [48:0] n1779_o;
  reg [5:0] n1830_o;
  reg n1854_o;
  wire [6:0] n1858_o;
  wire [6:0] n1859_o;
  wire [6:0] n1860_o;
  wire n1863_o;
  wire [5:0] n1865_o;
  wire [7:0] n1867_o;
  wire [5:0] n1868_o;
  wire [7:0] n1869_o;
  wire [5:0] n1870_o;
  wire n1880_o;
  wire [5:0] n1882_o;
  wire [5:0] n1883_o;
  wire int_b_n1884;
  wire int_b_n1886;
  wire int_b_n1887;
  wire int_b_n1888;
  wire int_b_tf_o;
  wire int_b_ext_int_o;
  wire int_b_tim_int_o;
  wire int_b_int_pending_o;
  wire int_b_int_in_progress_o;
  wire n1898_o;
  wire n1899_o;
  wire n1900_o;
  wire n1903_o;
  wire n1904_o;
  wire n1905_o;
  wire n1906_o;
  wire n1907_o;
  wire n1910_o;
  wire n1911_o;
  wire n1914_o;
  wire n1916_o;
  wire n1919_o;
  wire n1921_o;
  wire n1923_o;
  wire n1925_o;
  wire n1927_o;
  wire n1928_o;
  wire n1929_o;
  wire n1932_o;
  wire n1935_o;
  wire n1937_o;
  wire n1939_o;
  wire n1941_o;
  wire n1942_o;
  wire n1943_o;
  wire n1944_o;
  wire n1945_o;
  wire n1948_o;
  wire n1950_o;
  wire n1953_o;
  wire n1955_o;
  wire n1956_o;
  wire n1957_o;
  wire n1958_o;
  wire n1959_o;
  wire n1962_o;
  wire n1965_o;
  wire n1968_o;
  wire n1970_o;
  wire n1971_o;
  wire n1972_o;
  wire n1973_o;
  wire n1974_o;
  wire n1975_o;
  wire n1976_o;
  wire n1979_o;
  wire n1981_o;
  wire [4:0] n1982_o;
  reg n1984_o;
  reg n1987_o;
  reg n1990_o;
  reg n1993_o;
  reg n1996_o;
  reg n1999_o;
  reg n2002_o;
  reg n2005_o;
  reg n2008_o;
  wire n2015_o;
  wire n2016_o;
  wire n2018_o;
  wire n2019_o;
  wire n2020_o;
  wire [2:0] n2021_o;
  wire n2022_o;
  wire [2:0] n2024_o;
  wire [2:0] n2025_o;
  localparam [7:0] n2026_o = 8'b00000000;
  wire [4:0] n2027_o;
  wire n2030_o;
  wire [7:0] n2032_o;
  localparam [7:0] n2033_o = 8'bX;
  wire [7:0] n2034_o;
  wire n2038_o;
  wire n2040_o;
  wire n2041_o;
  wire n2043_o;
  wire n2050_o;
  wire n2053_o;
  wire [1:0] n2056_o;
  wire n2058_o;
  wire n2063_o;
  wire n2067_o;
  wire n2070_o;
  wire n2072_o;
  wire [2:0] n2073_o;
  reg n2076_o;
  reg n2079_o;
  reg n2082_o;
  reg n2083_o;
  reg n2086_o;
  reg [3:0] n2089_o;
  reg n2091_o;
  reg [1:0] n2093_o;
  reg n2095_o;
  reg n2098_o;
  reg n2101_o;
  wire n2103_o;
  wire n2105_o;
  wire n2109_o;
  wire n2112_o;
  wire n2114_o;
  wire [1:0] n2115_o;
  reg n2118_o;
  reg n2121_o;
  reg n2124_o;
  reg [3:0] n2127_o;
  reg n2129_o;
  reg n2131_o;
  reg n2134_o;
  reg n2137_o;
  wire n2139_o;
  wire n2141_o;
  wire n2143_o;
  wire [3:0] n2145_o;
  wire n2147_o;
  wire n2149_o;
  wire n2151_o;
  wire n2153_o;
  wire n2155_o;
  wire n2156_o;
  wire n2157_o;
  wire n2159_o;
  wire n2166_o;
  wire n2169_o;
  wire [1:0] n2172_o;
  wire n2174_o;
  wire n2179_o;
  wire n2184_o;
  wire [2:0] n2185_o;
  reg n2188_o;
  reg n2191_o;
  reg n2194_o;
  reg n2195_o;
  reg n2198_o;
  reg [3:0] n2201_o;
  reg [1:0] n2203_o;
  wire n2205_o;
  wire n2207_o;
  wire n2212_o;
  wire [1:0] n2213_o;
  reg n2216_o;
  reg n2219_o;
  reg n2222_o;
  reg [3:0] n2225_o;
  wire n2227_o;
  wire n2229_o;
  wire n2231_o;
  wire [3:0] n2233_o;
  wire n2235_o;
  wire n2236_o;
  wire n2238_o;
  wire [1:0] n2239_o;
  wire n2241_o;
  wire n2242_o;
  wire n2243_o;
  wire n2246_o;
  wire n2249_o;
  wire n2252_o;
  wire n2255_o;
  wire n2257_o;
  wire n2259_o;
  wire n2261_o;
  wire n2263_o;
  wire n2266_o;
  wire n2269_o;
  wire n2271_o;
  wire n2273_o;
  wire n2275_o;
  wire n2277_o;
  wire n2279_o;
  wire n2281_o;
  wire n2283_o;
  wire [1:0] n2284_o;
  wire n2286_o;
  wire n2287_o;
  wire n2288_o;
  wire n2291_o;
  wire n2294_o;
  wire n2297_o;
  wire n2299_o;
  wire n2301_o;
  wire n2303_o;
  wire [2:0] n2304_o;
  reg n2308_o;
  reg n2312_o;
  reg n2314_o;
  reg n2316_o;
  reg n2318_o;
  reg [3:0] n2321_o;
  wire n2323_o;
  wire n2325_o;
  wire n2327_o;
  wire n2329_o;
  wire n2331_o;
  wire n2333_o;
  wire n2335_o;
  wire n2337_o;
  wire [3:0] n2339_o;
  wire n2341_o;
  wire n2343_o;
  wire n2345_o;
  wire n2347_o;
  wire n2348_o;
  wire n2349_o;
  wire n2352_o;
  wire n2354_o;
  wire n2356_o;
  wire n2358_o;
  wire [2:0] n2359_o;
  reg n2362_o;
  reg n2365_o;
  reg n2368_o;
  reg n2371_o;
  reg n2374_o;
  reg [1:0] n2378_o;
  reg n2381_o;
  reg n2383_o;
  reg n2387_o;
  localparam [7:0] n2389_o = 8'b00000000;
  wire n2394_o;
  wire n2395_o;
  wire n2396_o;
  wire [4:0] n2397_o;
  wire n2399_o;
  wire [7:0] n2400_o;
  wire [7:0] n2401_o;
  wire n2403_o;
  wire n2405_o;
  wire n2406_o;
  wire [4:0] n2408_o;
  wire [2:0] n2409_o;
  wire [7:0] n2410_o;
  wire [7:0] n2412_o;
  wire n2415_o;
  wire n2417_o;
  wire [1:0] n2418_o;
  reg n2420_o;
  reg n2423_o;
  reg n2426_o;
  reg n2429_o;
  reg [7:0] n2430_o;
  reg n2432_o;
  reg n2434_o;
  wire n2436_o;
  wire n2437_o;
  wire n2439_o;
  wire n2441_o;
  wire n2443_o;
  wire n2445_o;
  wire n2447_o;
  wire n2449_o;
  wire [1:0] n2451_o;
  wire n2453_o;
  wire n2455_o;
  wire n2457_o;
  wire [7:0] n2458_o;
  wire n2459_o;
  wire n2461_o;
  wire n2463_o;
  wire n2465_o;
  wire n2467_o;
  wire n2470_o;
  wire n2473_o;
  wire [3:0] n2476_o;
  wire n2478_o;
  wire n2480_o;
  wire n2483_o;
  wire n2485_o;
  wire n2487_o;
  wire n2488_o;
  wire n2489_o;
  wire n2492_o;
  wire n2495_o;
  wire n2497_o;
  wire n2499_o;
  wire n2501_o;
  wire n2503_o;
  wire n2506_o;
  wire n2509_o;
  wire [3:0] n2512_o;
  wire n2514_o;
  wire n2516_o;
  wire n2517_o;
  wire n2519_o;
  wire n2522_o;
  wire n2524_o;
  wire n2526_o;
  wire n2527_o;
  wire n2528_o;
  wire n2529_o;
  wire n2531_o;
  wire n2534_o;
  wire n2537_o;
  wire n2539_o;
  wire n2541_o;
  wire n2543_o;
  wire n2545_o;
  wire n2547_o;
  wire n2548_o;
  wire n2551_o;
  wire n2554_o;
  wire n2556_o;
  wire [3:0] n2559_o;
  wire n2561_o;
  wire n2563_o;
  wire [2:0] n2564_o;
  reg n2567_o;
  reg n2569_o;
  reg n2572_o;
  reg [3:0] n2574_o;
  reg n2578_o;
  reg n2581_o;
  reg n2584_o;
  reg n2586_o;
  reg n2589_o;
  wire n2591_o;
  wire n2592_o;
  wire n2595_o;
  wire n2598_o;
  wire n2600_o;
  wire n2601_o;
  wire n2602_o;
  wire n2605_o;
  wire n2608_o;
  wire n2610_o;
  wire [1:0] n2611_o;
  reg n2613_o;
  reg n2615_o;
  reg n2618_o;
  reg n2620_o;
  reg [3:0] n2623_o;
  reg n2625_o;
  wire n2627_o;
  wire n2629_o;
  wire n2630_o;
  wire n2633_o;
  wire n2636_o;
  wire n2638_o;
  wire n2640_o;
  wire n2642_o;
  wire n2644_o;
  wire n2645_o;
  wire n2648_o;
  wire n2651_o;
  wire n2653_o;
  wire n2655_o;
  wire n2657_o;
  wire n2658_o;
  wire n2660_o;
  wire n2663_o;
  wire [1:0] n2664_o;
  reg n2667_o;
  reg n2670_o;
  reg n2673_o;
  reg [3:0] n2676_o;
  reg n2679_o;
  reg [3:0] n2682_o;
  wire n2683_o;
  reg n2684_o;
  reg n2687_o;
  wire n2689_o;
  wire n2690_o;
  wire n2696_o;
  wire n2699_o;
  wire n2701_o;
  wire n2703_o;
  wire n2705_o;
  wire n2707_o;
  wire [3:0] n2709_o;
  wire n2711_o;
  wire [3:0] n2713_o;
  wire n2714_o;
  wire n2715_o;
  wire n2717_o;
  wire n2719_o;
  wire n2721_o;
  wire n2723_o;
  wire n2724_o;
  wire n2725_o;
  wire n2728_o;
  wire n2731_o;
  wire n2733_o;
  wire n2735_o;
  wire n2737_o;
  wire n2739_o;
  wire n2742_o;
  wire n2744_o;
  wire n2746_o;
  wire n2747_o;
  wire n2748_o;
  wire n2749_o;
  wire n2752_o;
  wire n2755_o;
  wire n2758_o;
  wire n2760_o;
  wire n2762_o;
  wire n2764_o;
  wire n2766_o;
  wire n2769_o;
  wire n2772_o;
  wire n2774_o;
  wire n2776_o;
  wire n2777_o;
  wire n2780_o;
  wire n2783_o;
  wire n2785_o;
  wire n2786_o;
  wire n2787_o;
  wire n2789_o;
  wire n2796_o;
  wire n2799_o;
  wire [1:0] n2802_o;
  wire n2804_o;
  wire [1:0] n2805_o;
  wire n2807_o;
  wire n2810_o;
  wire n2813_o;
  wire n2815_o;
  wire [1:0] n2816_o;
  wire n2818_o;
  wire n2821_o;
  wire n2824_o;
  wire n2826_o;
  wire [2:0] n2827_o;
  reg n2829_o;
  reg n2831_o;
  reg n2834_o;
  reg n2835_o;
  reg n2837_o;
  reg [3:0] n2840_o;
  reg [1:0] n2842_o;
  reg n2844_o;
  wire n2846_o;
  wire n2847_o;
  wire n2849_o;
  wire n2852_o;
  wire n2855_o;
  wire n2857_o;
  wire n2858_o;
  wire n2864_o;
  wire n2867_o;
  wire n2869_o;
  wire n2871_o;
  wire n2873_o;
  wire n2875_o;
  wire n2877_o;
  wire n2878_o;
  wire n2880_o;
  wire n2881_o;
  wire n2884_o;
  wire n2885_o;
  wire n2886_o;
  wire n2888_o;
  wire n2889_o;
  wire n2895_o;
  wire n2898_o;
  wire n2900_o;
  wire n2902_o;
  wire n2904_o;
  wire n2906_o;
  wire n2908_o;
  wire n2909_o;
  wire n2911_o;
  wire n2912_o;
  wire [3:0] n2915_o;
  wire n2918_o;
  wire [3:0] n2920_o;
  wire n2922_o;
  wire n2923_o;
  wire n2929_o;
  wire n2932_o;
  wire n2934_o;
  wire n2936_o;
  wire [3:0] n2938_o;
  wire n2940_o;
  wire n2942_o;
  wire n2944_o;
  wire [4:0] n2946_o;
  wire [2:0] n2947_o;
  wire [7:0] n2948_o;
  wire n2950_o;
  wire [1:0] n2951_o;
  reg n2954_o;
  reg n2957_o;
  reg n2960_o;
  reg [7:0] n2961_o;
  reg n2963_o;
  wire n2965_o;
  wire n2967_o;
  wire n2969_o;
  wire [7:0] n2970_o;
  wire n2971_o;
  wire n2973_o;
  wire n2974_o;
  wire n2976_o;
  wire n2979_o;
  wire [1:0] n2982_o;
  wire n2984_o;
  wire n2987_o;
  wire n2990_o;
  wire n2992_o;
  wire n2994_o;
  wire [1:0] n2996_o;
  wire n2998_o;
  wire n3000_o;
  wire n3001_o;
  wire n3003_o;
  wire n3006_o;
  wire n3008_o;
  wire n3009_o;
  wire n3015_o;
  wire n3018_o;
  wire n3020_o;
  wire n3022_o;
  wire n3024_o;
  wire n3026_o;
  wire n3027_o;
  wire n3029_o;
  wire n3032_o;
  wire n3034_o;
  wire n3035_o;
  wire n3041_o;
  wire n3044_o;
  wire n3046_o;
  wire n3048_o;
  wire n3050_o;
  wire n3052_o;
  wire n3053_o;
  wire n3055_o;
  wire n3058_o;
  wire n3060_o;
  wire n3061_o;
  wire n3067_o;
  wire n3070_o;
  wire n3072_o;
  wire n3074_o;
  wire n3076_o;
  wire n3078_o;
  wire n3079_o;
  wire n3080_o;
  wire [3:0] n3083_o;
  wire n3084_o;
  wire n3086_o;
  wire n3087_o;
  wire n3090_o;
  wire n3091_o;
  wire n3092_o;
  wire n3094_o;
  wire n3095_o;
  wire n3101_o;
  wire n3104_o;
  wire n3106_o;
  wire n3108_o;
  wire n3110_o;
  wire n3112_o;
  wire n3114_o;
  wire n3115_o;
  wire n3117_o;
  wire n3120_o;
  wire n3123_o;
  wire n3125_o;
  wire n3126_o;
  wire n3132_o;
  wire n3135_o;
  wire n3137_o;
  wire n3139_o;
  wire n3141_o;
  wire n3143_o;
  wire n3145_o;
  wire n3146_o;
  wire n3148_o;
  wire n3149_o;
  wire n3152_o;
  wire n3155_o;
  wire n3156_o;
  wire n3157_o;
  wire n3159_o;
  wire n3160_o;
  wire n3166_o;
  wire n3169_o;
  wire n3171_o;
  wire n3173_o;
  wire n3175_o;
  wire n3177_o;
  wire n3179_o;
  wire n3181_o;
  wire n3183_o;
  wire n3184_o;
  wire n3187_o;
  wire n3189_o;
  wire n3190_o;
  wire n3191_o;
  wire n3193_o;
  wire n3200_o;
  wire n3203_o;
  wire [1:0] n3206_o;
  wire n3208_o;
  wire n3213_o;
  wire [1:0] n3214_o;
  reg n3217_o;
  reg n3220_o;
  reg n3221_o;
  reg n3224_o;
  reg [1:0] n3226_o;
  wire n3228_o;
  wire n3230_o;
  wire n3233_o;
  wire n3236_o;
  wire n3239_o;
  wire n3241_o;
  wire n3243_o;
  wire n3246_o;
  wire n3249_o;
  wire n3252_o;
  wire n3254_o;
  wire n3255_o;
  wire n3256_o;
  wire n3258_o;
  wire n3265_o;
  wire n3268_o;
  wire [1:0] n3271_o;
  wire n3273_o;
  wire n3275_o;
  wire [1:0] n3276_o;
  reg n3279_o;
  reg n3280_o;
  reg n3282_o;
  reg [1:0] n3284_o;
  reg n3287_o;
  wire n3289_o;
  wire n3290_o;
  wire n3292_o;
  wire n3293_o;
  wire n3294_o;
  wire n3295_o;
  wire n3297_o;
  wire n3304_o;
  wire n3307_o;
  wire [1:0] n3310_o;
  wire n3311_o;
  wire n3313_o;
  wire [1:0] n3315_o;
  wire n3317_o;
  wire n3318_o;
  wire n3321_o;
  wire n3323_o;
  wire n3325_o;
  wire n3328_o;
  wire n3331_o;
  wire n3333_o;
  wire n3335_o;
  wire n3336_o;
  wire n3339_o;
  wire n3342_o;
  wire n3345_o;
  wire n3348_o;
  wire n3350_o;
  wire n3352_o;
  wire n3354_o;
  wire n3356_o;
  wire n3358_o;
  wire n3359_o;
  wire [1:0] n3361_o;
  wire [3:0] n3362_o;
  wire n3365_o;
  wire n3368_o;
  wire n3371_o;
  wire [2:0] n3372_o;
  wire [1:0] n3373_o;
  wire [1:0] n3374_o;
  wire [1:0] n3375_o;
  reg [1:0] n3376_o;
  wire n3378_o;
  wire n3380_o;
  wire n3382_o;
  wire [2:0] n3383_o;
  reg n3386_o;
  reg n3390_o;
  wire [1:0] n3391_o;
  wire [1:0] n3392_o;
  wire [1:0] n3393_o;
  reg [1:0] n3394_o;
  wire [1:0] n3395_o;
  wire [1:0] n3396_o;
  wire [1:0] n3397_o;
  reg [1:0] n3398_o;
  wire [3:0] n3399_o;
  wire [3:0] n3400_o;
  wire [3:0] n3401_o;
  reg [3:0] n3402_o;
  reg n3404_o;
  reg n3408_o;
  wire n3410_o;
  wire n3412_o;
  wire n3413_o;
  wire n3416_o;
  wire n3418_o;
  wire n3420_o;
  wire [7:0] n3421_o;
  wire [7:0] n3422_o;
  wire n3423_o;
  wire n3424_o;
  wire n3426_o;
  wire n3427_o;
  wire [1:0] n3428_o;
  wire [7:0] n3430_o;
  wire n3432_o;
  wire n3435_o;
  wire n3437_o;
  wire [2:0] n3438_o;
  reg n3442_o;
  wire [3:0] n3443_o;
  wire [3:0] n3444_o;
  wire [3:0] n3445_o;
  wire [3:0] n3446_o;
  reg [3:0] n3447_o;
  wire [3:0] n3448_o;
  wire [3:0] n3449_o;
  wire [3:0] n3450_o;
  wire [3:0] n3451_o;
  reg [3:0] n3452_o;
  reg n3455_o;
  reg n3459_o;
  wire n3461_o;
  wire n3463_o;
  wire [1:0] n3464_o;
  reg n3467_o;
  reg n3470_o;
  reg n3473_o;
  reg n3477_o;
  wire n3479_o;
  wire n3481_o;
  wire n3483_o;
  wire n3485_o;
  wire [7:0] n3486_o;
  wire [7:0] n3487_o;
  wire n3488_o;
  wire n3489_o;
  wire n3491_o;
  wire n3492_o;
  wire n3494_o;
  wire n3495_o;
  wire n3496_o;
  wire [1:0] n3499_o;
  wire n3502_o;
  wire [1:0] n3504_o;
  wire n3506_o;
  wire n3509_o;
  wire n3512_o;
  wire n3514_o;
  wire n3516_o;
  wire [1:0] n3518_o;
  wire n3520_o;
  wire n3522_o;
  wire n3523_o;
  wire n3524_o;
  wire n3527_o;
  wire n3530_o;
  wire n3531_o;
  wire n3533_o;
  wire n3534_o;
  wire n3537_o;
  wire n3540_o;
  wire n3542_o;
  wire [1:0] n3543_o;
  reg n3545_o;
  reg n3548_o;
  reg n3551_o;
  wire n3553_o;
  wire n3554_o;
  wire n3555_o;
  wire n3558_o;
  wire n3561_o;
  wire n3564_o;
  wire n3567_o;
  wire n3569_o;
  wire n3571_o;
  wire n3573_o;
  wire n3575_o;
  wire n3577_o;
  wire n3578_o;
  wire n3579_o;
  wire n3581_o;
  wire n3583_o;
  wire n3586_o;
  wire n3588_o;
  wire n3590_o;
  wire n3591_o;
  wire n3592_o;
  wire n3594_o;
  wire n3601_o;
  wire n3604_o;
  wire [1:0] n3607_o;
  wire n3609_o;
  wire n3614_o;
  wire n3619_o;
  wire [2:0] n3620_o;
  reg n3623_o;
  reg n3626_o;
  reg n3629_o;
  reg n3630_o;
  reg n3633_o;
  reg [3:0] n3636_o;
  reg [1:0] n3638_o;
  wire n3640_o;
  wire n3642_o;
  wire n3647_o;
  wire [1:0] n3648_o;
  reg n3651_o;
  reg n3654_o;
  reg n3657_o;
  reg [3:0] n3660_o;
  wire n3662_o;
  wire n3664_o;
  wire n3666_o;
  wire [3:0] n3668_o;
  wire n3670_o;
  wire n3671_o;
  wire n3673_o;
  wire [1:0] n3674_o;
  wire n3676_o;
  wire n3677_o;
  wire n3678_o;
  wire n3681_o;
  wire n3684_o;
  wire n3687_o;
  wire n3690_o;
  wire n3692_o;
  wire n3694_o;
  wire n3696_o;
  wire n3698_o;
  wire n3701_o;
  wire n3704_o;
  wire n3706_o;
  wire n3708_o;
  wire n3710_o;
  wire n3712_o;
  wire n3714_o;
  wire n3716_o;
  wire n3718_o;
  wire [1:0] n3719_o;
  wire n3721_o;
  wire n3722_o;
  wire n3723_o;
  wire n3726_o;
  wire n3729_o;
  wire n3732_o;
  wire n3734_o;
  wire n3736_o;
  wire n3738_o;
  wire [2:0] n3739_o;
  reg n3743_o;
  reg n3747_o;
  reg n3749_o;
  reg n3751_o;
  reg n3753_o;
  reg [3:0] n3756_o;
  wire n3758_o;
  wire n3760_o;
  wire n3762_o;
  wire n3764_o;
  wire n3766_o;
  wire n3768_o;
  wire n3770_o;
  wire n3772_o;
  wire [3:0] n3774_o;
  wire n3776_o;
  wire n3778_o;
  wire n3780_o;
  wire n3782_o;
  wire n3784_o;
  wire n3787_o;
  wire n3790_o;
  wire n3792_o;
  wire n3793_o;
  wire n3794_o;
  wire n3797_o;
  wire n3798_o;
  wire n3800_o;
  wire n3801_o;
  wire n3802_o;
  wire n3803_o;
  wire n3804_o;
  wire n3807_o;
  wire n3810_o;
  wire n3813_o;
  wire n3815_o;
  wire n3817_o;
  wire n3820_o;
  wire n3822_o;
  wire n3824_o;
  wire n3826_o;
  wire n3828_o;
  wire n3829_o;
  wire n3831_o;
  wire n3833_o;
  wire n3835_o;
  wire [2:0] n3836_o;
  reg n3839_o;
  reg n3842_o;
  reg n3845_o;
  reg n3848_o;
  reg [1:0] n3852_o;
  reg n3855_o;
  wire n3856_o;
  wire n3859_o;
  wire n3862_o;
  wire n3864_o;
  wire n3866_o;
  wire [1:0] n3867_o;
  reg n3870_o;
  reg n3873_o;
  reg n3875_o;
  reg n3878_o;
  reg n3880_o;
  wire n3881_o;
  wire n3882_o;
  wire n3884_o;
  wire n3886_o;
  wire n3888_o;
  wire n3890_o;
  wire [1:0] n3892_o;
  wire n3894_o;
  wire n3896_o;
  wire n3898_o;
  wire n3900_o;
  wire n3902_o;
  wire n3903_o;
  wire n3906_o;
  wire n3908_o;
  wire n3911_o;
  wire n3914_o;
  wire n3917_o;
  wire [3:0] n3920_o;
  wire n3922_o;
  wire n3924_o;
  wire n3926_o;
  wire n3928_o;
  wire n3930_o;
  wire n3931_o;
  wire n3932_o;
  wire n3935_o;
  wire n3937_o;
  wire n3940_o;
  wire n3943_o;
  wire n3946_o;
  wire [3:0] n3949_o;
  wire n3951_o;
  wire n3953_o;
  wire n3955_o;
  wire n3957_o;
  wire n3959_o;
  wire n3960_o;
  wire n3963_o;
  wire n3966_o;
  wire n3968_o;
  wire n3970_o;
  wire n3972_o;
  wire n3974_o;
  wire n3975_o;
  wire n3977_o;
  wire n3980_o;
  wire n3982_o;
  wire n3984_o;
  wire n3987_o;
  wire n3989_o;
  wire n3991_o;
  wire n3992_o;
  wire n3995_o;
  wire n3998_o;
  wire n4000_o;
  wire n4002_o;
  wire n4004_o;
  wire n4006_o;
  wire n4009_o;
  wire n4012_o;
  wire n4014_o;
  wire n4015_o;
  wire n4016_o;
  wire n4018_o;
  wire n4025_o;
  wire n4028_o;
  wire [1:0] n4031_o;
  wire n4033_o;
  wire n4034_o;
  wire n4037_o;
  wire n4039_o;
  wire n4040_o;
  wire [3:0] n4043_o;
  wire n4045_o;
  wire [2:0] n4046_o;
  reg n4049_o;
  reg n4052_o;
  reg n4055_o;
  reg n4056_o;
  reg n4059_o;
  reg [3:0] n4061_o;
  reg n4063_o;
  reg [1:0] n4065_o;
  reg n4068_o;
  wire n4070_o;
  wire n4071_o;
  wire n4072_o;
  wire n4074_o;
  wire n4081_o;
  wire n4084_o;
  wire [1:0] n4087_o;
  wire n4089_o;
  wire n4094_o;
  wire n4099_o;
  wire [2:0] n4100_o;
  reg n4103_o;
  reg n4106_o;
  reg n4109_o;
  reg n4110_o;
  reg n4113_o;
  reg [3:0] n4116_o;
  reg [1:0] n4118_o;
  wire n4120_o;
  wire n4122_o;
  wire n4127_o;
  wire [1:0] n4128_o;
  reg n4131_o;
  reg n4134_o;
  reg n4137_o;
  reg [3:0] n4140_o;
  wire n4142_o;
  wire n4144_o;
  wire n4146_o;
  wire [3:0] n4148_o;
  wire n4150_o;
  wire [62:0] n4151_o;
  reg n4153_o;
  reg n4156_o;
  reg n4159_o;
  reg n4162_o;
  reg n4165_o;
  reg n4168_o;
  reg n4171_o;
  reg n4174_o;
  reg n4177_o;
  reg n4179_o;
  reg n4181_o;
  reg n4184_o;
  reg n4187_o;
  reg n4190_o;
  reg n4193_o;
  reg n4196_o;
  reg n4199_o;
  reg n4202_o;
  reg n4205_o;
  reg n4208_o;
  reg n4211_o;
  reg n4214_o;
  reg n4217_o;
  reg n4220_o;
  reg n4223_o;
  reg [3:0] n4227_o;
  reg n4230_o;
  reg n4233_o;
  reg n4236_o;
  reg n4239_o;
  reg n4242_o;
  reg n4246_o;
  reg n4251_o;
  reg n4255_o;
  reg n4258_o;
  reg n4261_o;
  reg [3:0] n4271_o;
  wire n4273_o;
  reg n4274_o;
  wire [1:0] n4275_o;
  reg [1:0] n4277_o;
  reg n4280_o;
  reg n4283_o;
  reg [1:0] n4286_o;
  reg n4289_o;
  reg n4292_o;
  reg n4295_o;
  reg n4298_o;
  reg n4301_o;
  reg n4304_o;
  reg n4307_o;
  reg n4310_o;
  reg n4313_o;
  reg n4316_o;
  reg n4319_o;
  reg n4322_o;
  reg n4347_o;
  reg n4350_o;
  reg n4353_o;
  reg n4356_o;
  reg n4359_o;
  reg n4362_o;
  reg n4365_o;
  reg n4368_o;
  reg n4371_o;
  reg [7:0] n4373_o;
  reg n4374_o;
  reg n4376_o;
  reg n4379_o;
  reg n4382_o;
  reg n4385_o;
  reg n4388_o;
  reg n4391_o;
  reg n4394_o;
  reg n4397_o;
  reg n4400_o;
  reg n4403_o;
  reg n4406_o;
  wire n4410_o;
  wire n4413_o;
  wire n4415_o;
  wire n4417_o;
  wire n4419_o;
  wire n4421_o;
  wire n4422_o;
  wire n4423_o;
  wire n4425_o;
  wire n4427_o;
  wire n4429_o;
  wire n4433_o;
  wire n4435_o;
  wire [7:0] n4449_o;
  wire n4451_o;
  wire n4452_o;
  wire n4453_o;
  wire n4454_o;
  wire [7:0] n4455_o;
  reg [7:0] n4456_q;
  wire n4457_o;
  reg n4458_q;
  reg n4459_q;
  wire n4460_o;
  reg n4461_q;
  wire n4462_o;
  reg n4463_q;
  wire [5:0] n4464_o;
  reg [5:0] n4465_q;
  wire [2:0] n4466_o;
  assign t0_dir_o = t0_dir_q;
  assign data_o = n4449_o;
  assign alu_write_accu_o = n4153_o;
  assign alu_write_shadow_o = n4156_o;
  assign alu_write_temp_reg_o = n4159_o;
  assign alu_read_alu_o = n4162_o;
  assign bus_write_bus_o = n4165_o;
  assign bus_read_bus_o = n4454_o;
  assign bus_ibf_int_o = n4168_o;
  assign bus_en_dma_o = n4171_o;
  assign bus_en_flags_o = n4174_o;
  assign bus_write_sts_o = n4177_o;
  assign dm_write_dmem_addr_o = n4179_o;
  assign dm_write_dmem_o = n4451_o;
  assign dm_read_dmem_o = n4181_o;
  assign p1_write_p1_o = n4184_o;
  assign p1_read_p1_o = n4187_o;
  assign p2_write_p2_o = n4190_o;
  assign p2_write_exp_o = n4193_o;
  assign p2_read_p2_o = n4196_o;
  assign p2_read_exp_o = n4199_o;
  assign pm_write_pcl_o = n4202_o;
  assign pm_read_pcl_o = n4205_o;
  assign pm_write_pch_o = n4208_o;
  assign pm_read_pch_o = n4211_o;
  assign pm_read_pmem_o = n1984_o;
  assign psw_read_psw_o = n4214_o;
  assign psw_read_sp_o = n4217_o;
  assign psw_write_psw_o = n4220_o;
  assign psw_write_sp_o = n4223_o;
  assign alu_op_o = n4227_o;
  assign alu_use_carry_o = n4230_o;
  assign alu_da_high_o = n4233_o;
  assign alu_accu_low_o = n4236_o;
  assign alu_p06_temp_reg_o = n4239_o;
  assign alu_p60_temp_reg_o = n4242_o;
  assign bus_output_pcl_o = n1987_o;
  assign bus_bidir_bus_o = n4246_o;
  assign clk_multi_cycle_o = opc_multi_cycle_s;
  assign clk_assert_psen_o = n1990_o;
  assign clk_assert_prog_o = n4251_o;
  assign clk_assert_rd_o = n4255_o;
  assign clk_assert_wr_o = n4258_o;
  assign cnd_compute_take_o = n4261_o;
  assign cnd_branch_cond_o = n4271_o;
  assign cnd_comp_value_o = n4466_o;
  assign cnd_f1_o = f1_q;
  assign cnd_tf_o = tf_s;
  assign dm_addr_type_o = n4277_o;
  assign p1_read_reg_o = n4280_o;
  assign p2_read_reg_o = n4283_o;
  assign p2_output_pch_o = n1993_o;
  assign pm_inc_pc_o = n4452_o;
  assign pm_write_pmem_addr_o = n4453_o;
  assign pm_addr_type_o = n4286_o;
  assign psw_special_data_o = n4289_o;
  assign psw_inc_stackp_o = n4292_o;
  assign psw_dec_stackp_o = n4295_o;
  assign psw_write_carry_o = n4298_o;
  assign psw_write_aux_carry_o = n4301_o;
  assign psw_write_f0_o = n4304_o;
  assign psw_write_bs_o = n4307_o;
  assign tim_read_timer_o = n4310_o;
  assign tim_write_timer_o = n4313_o;
  assign tim_start_t_o = n4316_o;
  assign tim_start_cnt_o = n4319_o;
  assign tim_stop_tcnt_o = n4322_o;
  /* decoder.vhd:187:10  */
  assign opc_multi_cycle_s = n1880_o; // (signal)
  /* decoder.vhd:188:10  */
  assign opc_read_bus_s = n1996_o; // (signal)
  /* decoder.vhd:189:10  */
  assign opc_inj_int_s = n1999_o; // (signal)
  /* decoder.vhd:190:10  */
  assign opc_opcode_q = n4456_q; // (signal)
  /* decoder.vhd:191:10  */
  assign opc_mnemonic_s = n1882_o; // (signal)
  /* decoder.vhd:192:10  */
  assign last_cycle_s = n1900_o; // (signal)
  /* decoder.vhd:195:10  */
  assign assert_psen_s = n4347_o; // (signal)
  /* decoder.vhd:198:10  */
  assign branch_taken_s = n4350_o; // (signal)
  /* decoder.vhd:199:10  */
  assign branch_taken_q = n4458_q; // (signal)
  /* decoder.vhd:200:10  */
  assign pm_inc_pc_s = n2002_o; // (signal)
  /* decoder.vhd:201:10  */
  assign pm_write_pmem_addr_s = n2005_o; // (signal)
  /* decoder.vhd:203:10  */
  assign add_inc_pc_s = n4353_o; // (signal)
  /* decoder.vhd:205:10  */
  assign add_write_pmem_addr_s = n4356_o; // (signal)
  /* decoder.vhd:208:10  */
  assign clear_f1_s = n4359_o; // (signal)
  /* decoder.vhd:209:10  */
  assign cpl_f1_s = n4362_o; // (signal)
  /* decoder.vhd:210:10  */
  assign f1_q = n4459_q; // (signal)
  /* decoder.vhd:212:10  */
  assign clear_mb_s = n4365_o; // (signal)
  /* decoder.vhd:213:10  */
  assign set_mb_s = n4368_o; // (signal)
  /* decoder.vhd:214:10  */
  assign mb_q = n4461_q; // (signal)
  /* decoder.vhd:217:10  */
  assign ent0_clk_s = n4371_o; // (signal)
  /* decoder.vhd:218:10  */
  assign t0_dir_q = n4463_q; // (signal)
  /* decoder.vhd:220:10  */
  assign data_s = n4373_o; // (signal)
  /* decoder.vhd:221:10  */
  assign read_dec_s = n4374_o; // (signal)
  /* decoder.vhd:223:10  */
  assign tf_s = int_b_n1884; // (signal)
  /* decoder.vhd:225:10  */
  assign bus_read_bus_s = n2008_o; // (signal)
  /* decoder.vhd:226:10  */
  assign add_read_bus_s = n4376_o; // (signal)
  /* decoder.vhd:228:10  */
  assign dm_write_dmem_s = n4379_o; // (signal)
  /* decoder.vhd:230:10  */
  assign p2_output_exp_s = n4382_o; // (signal)
  /* decoder.vhd:232:10  */
  assign movx_first_cycle_s = n4385_o; // (signal)
  /* decoder.vhd:235:10  */
  assign jtf_executed_s = n4388_o; // (signal)
  /* decoder.vhd:236:10  */
  assign en_tcnti_s = n4391_o; // (signal)
  /* decoder.vhd:237:10  */
  assign dis_tcnti_s = n4394_o; // (signal)
  /* decoder.vhd:238:10  */
  assign en_i_s = n4397_o; // (signal)
  /* decoder.vhd:239:10  */
  assign dis_i_s = n4400_o; // (signal)
  /* decoder.vhd:240:10  */
  assign tim_int_s = int_b_n1886; // (signal)
  /* decoder.vhd:241:10  */
  assign retr_executed_s = n4403_o; // (signal)
  /* decoder.vhd:242:10  */
  assign int_executed_s = n4406_o; // (signal)
  /* decoder.vhd:243:10  */
  assign int_pending_s = int_b_n1887; // (signal)
  /* decoder.vhd:244:10  */
  assign int_in_progress_s = int_b_n1888; // (signal)
  /* decoder.vhd:247:10  */
  assign mnemonic_rec_s = n1860_o; // (signal)
  /* decoder.vhd:248:10  */
  assign mnemonic_q = n4465_q; // (signal)
  /* decoder_pack-p.vhd:419:7  */
  assign n1116_o = opc_opcode_q == 8'b10011000;
  /* decoder_pack-p.vhd:419:23  */
  assign n1118_o = opc_opcode_q == 8'b10011001;
  /* decoder_pack-p.vhd:419:23  */
  assign n1119_o = n1116_o | n1118_o;
  /* decoder_pack-p.vhd:420:23  */
  assign n1121_o = opc_opcode_q == 8'b10011010;
  /* decoder_pack-p.vhd:420:23  */
  assign n1122_o = n1119_o | n1121_o;
  /* decoder_pack-p.vhd:425:7  */
  assign n1124_o = opc_opcode_q == 8'b01110101;
  /* decoder_pack-p.vhd:429:7  */
  assign n1126_o = opc_opcode_q == 8'b00001000;
  /* decoder_pack-p.vhd:434:7  */
  assign n1128_o = opc_opcode_q == 8'b10000110;
  /* decoder_pack-p.vhd:439:7  */
  assign n1130_o = opc_opcode_q == 8'b10000000;
  /* decoder_pack-p.vhd:439:23  */
  assign n1132_o = opc_opcode_q == 8'b10000001;
  /* decoder_pack-p.vhd:439:23  */
  assign n1133_o = n1130_o | n1132_o;
  /* decoder_pack-p.vhd:439:36  */
  assign n1135_o = opc_opcode_q == 8'b10010000;
  /* decoder_pack-p.vhd:439:36  */
  assign n1136_o = n1133_o | n1135_o;
  /* decoder_pack-p.vhd:440:23  */
  assign n1138_o = opc_opcode_q == 8'b10010001;
  /* decoder_pack-p.vhd:440:23  */
  assign n1139_o = n1136_o | n1138_o;
  /* decoder_pack-p.vhd:445:7  */
  assign n1141_o = opc_opcode_q == 8'b10001000;
  /* decoder_pack-p.vhd:445:23  */
  assign n1143_o = opc_opcode_q == 8'b10001001;
  /* decoder_pack-p.vhd:445:23  */
  assign n1144_o = n1141_o | n1143_o;
  /* decoder_pack-p.vhd:446:23  */
  assign n1146_o = opc_opcode_q == 8'b10001010;
  /* decoder_pack-p.vhd:446:23  */
  assign n1147_o = n1144_o | n1146_o;
  /* decoder_pack-p.vhd:451:7  */
  assign n1149_o = opc_opcode_q == 8'b00111001;
  /* decoder_pack-p.vhd:451:23  */
  assign n1151_o = opc_opcode_q == 8'b00111010;
  /* decoder_pack-p.vhd:451:23  */
  assign n1152_o = n1149_o | n1151_o;
  /* decoder_pack-p.vhd:451:36  */
  assign n1154_o = opc_opcode_q == 8'b00000010;
  /* decoder_pack-p.vhd:451:36  */
  assign n1155_o = n1152_o | n1154_o;
  /* decoder_pack-p.vhd:457:7  */
  assign n1157_o = opc_opcode_q == 8'b11100101;
  /* decoder_pack-p.vhd:457:23  */
  assign n1159_o = opc_opcode_q == 8'b11110101;
  /* decoder_pack-p.vhd:457:23  */
  assign n1160_o = n1157_o | n1159_o;
  assign n1161_o = {n1160_o, n1155_o, n1147_o, n1139_o, n1128_o, n1126_o, n1124_o, n1122_o};
  /* decoder_pack-p.vhd:417:5  */
  always @*
    case (n1161_o)
      8'b10000000: n1171_o = 6'b110010;
      8'b01000000: n1171_o = 6'b101110;
      8'b00100000: n1171_o = 6'b101100;
      8'b00010000: n1171_o = 6'b101000;
      8'b00001000: n1171_o = 6'b011011;
      8'b00000100: n1171_o = 6'b010101;
      8'b00000010: n1171_o = 6'b010010;
      8'b00000001: n1171_o = 6'b000101;
      default: n1171_o = 6'b000000;
    endcase
  /* decoder_pack-p.vhd:417:5  */
  always @*
    case (n1161_o)
      8'b10000000: n1180_o = 1'b0;
      8'b01000000: n1180_o = 1'b1;
      8'b00100000: n1180_o = 1'b1;
      8'b00010000: n1180_o = 1'b1;
      8'b00001000: n1180_o = 1'b1;
      8'b00000100: n1180_o = 1'b1;
      8'b00000010: n1180_o = 1'b0;
      8'b00000001: n1180_o = 1'b1;
      default: n1180_o = 1'b0;
    endcase
  /* decoder_pack-p.vhd:466:19  */
  assign n1183_o = n1171_o == 6'b000000;
  /* decoder_pack-p.vhd:123:7  */
  assign n1193_o = opc_opcode_q == 8'b01101000;
  /* decoder_pack-p.vhd:123:23  */
  assign n1195_o = opc_opcode_q == 8'b01101001;
  /* decoder_pack-p.vhd:123:23  */
  assign n1196_o = n1193_o | n1195_o;
  /* decoder_pack-p.vhd:123:36  */
  assign n1198_o = opc_opcode_q == 8'b01101010;
  /* decoder_pack-p.vhd:123:36  */
  assign n1199_o = n1196_o | n1198_o;
  /* decoder_pack-p.vhd:123:49  */
  assign n1201_o = opc_opcode_q == 8'b01101011;
  /* decoder_pack-p.vhd:123:49  */
  assign n1202_o = n1199_o | n1201_o;
  /* decoder_pack-p.vhd:123:62  */
  assign n1204_o = opc_opcode_q == 8'b01101100;
  /* decoder_pack-p.vhd:123:62  */
  assign n1205_o = n1202_o | n1204_o;
  /* decoder_pack-p.vhd:124:23  */
  assign n1207_o = opc_opcode_q == 8'b01101101;
  /* decoder_pack-p.vhd:124:23  */
  assign n1208_o = n1205_o | n1207_o;
  /* decoder_pack-p.vhd:124:36  */
  assign n1210_o = opc_opcode_q == 8'b01101110;
  /* decoder_pack-p.vhd:124:36  */
  assign n1211_o = n1208_o | n1210_o;
  /* decoder_pack-p.vhd:124:49  */
  assign n1213_o = opc_opcode_q == 8'b01101111;
  /* decoder_pack-p.vhd:124:49  */
  assign n1214_o = n1211_o | n1213_o;
  /* decoder_pack-p.vhd:124:62  */
  assign n1216_o = opc_opcode_q == 8'b01100000;
  /* decoder_pack-p.vhd:124:62  */
  assign n1217_o = n1214_o | n1216_o;
  /* decoder_pack-p.vhd:125:23  */
  assign n1219_o = opc_opcode_q == 8'b01100001;
  /* decoder_pack-p.vhd:125:23  */
  assign n1220_o = n1217_o | n1219_o;
  /* decoder_pack-p.vhd:125:36  */
  assign n1222_o = opc_opcode_q == 8'b01111000;
  /* decoder_pack-p.vhd:125:36  */
  assign n1223_o = n1220_o | n1222_o;
  /* decoder_pack-p.vhd:126:23  */
  assign n1225_o = opc_opcode_q == 8'b01111001;
  /* decoder_pack-p.vhd:126:23  */
  assign n1226_o = n1223_o | n1225_o;
  /* decoder_pack-p.vhd:126:36  */
  assign n1228_o = opc_opcode_q == 8'b01111010;
  /* decoder_pack-p.vhd:126:36  */
  assign n1229_o = n1226_o | n1228_o;
  /* decoder_pack-p.vhd:126:49  */
  assign n1231_o = opc_opcode_q == 8'b01111011;
  /* decoder_pack-p.vhd:126:49  */
  assign n1232_o = n1229_o | n1231_o;
  /* decoder_pack-p.vhd:126:62  */
  assign n1234_o = opc_opcode_q == 8'b01111100;
  /* decoder_pack-p.vhd:126:62  */
  assign n1235_o = n1232_o | n1234_o;
  /* decoder_pack-p.vhd:127:23  */
  assign n1237_o = opc_opcode_q == 8'b01111101;
  /* decoder_pack-p.vhd:127:23  */
  assign n1238_o = n1235_o | n1237_o;
  /* decoder_pack-p.vhd:127:36  */
  assign n1240_o = opc_opcode_q == 8'b01111110;
  /* decoder_pack-p.vhd:127:36  */
  assign n1241_o = n1238_o | n1240_o;
  /* decoder_pack-p.vhd:127:49  */
  assign n1243_o = opc_opcode_q == 8'b01111111;
  /* decoder_pack-p.vhd:127:49  */
  assign n1244_o = n1241_o | n1243_o;
  /* decoder_pack-p.vhd:127:62  */
  assign n1246_o = opc_opcode_q == 8'b01110000;
  /* decoder_pack-p.vhd:127:62  */
  assign n1247_o = n1244_o | n1246_o;
  /* decoder_pack-p.vhd:128:23  */
  assign n1249_o = opc_opcode_q == 8'b01110001;
  /* decoder_pack-p.vhd:128:23  */
  assign n1250_o = n1247_o | n1249_o;
  /* decoder_pack-p.vhd:132:7  */
  assign n1252_o = opc_opcode_q == 8'b00000011;
  /* decoder_pack-p.vhd:132:23  */
  assign n1254_o = opc_opcode_q == 8'b00010011;
  /* decoder_pack-p.vhd:132:23  */
  assign n1255_o = n1252_o | n1254_o;
  /* decoder_pack-p.vhd:138:7  */
  assign n1257_o = opc_opcode_q == 8'b01011000;
  /* decoder_pack-p.vhd:138:23  */
  assign n1259_o = opc_opcode_q == 8'b01011001;
  /* decoder_pack-p.vhd:138:23  */
  assign n1260_o = n1257_o | n1259_o;
  /* decoder_pack-p.vhd:138:36  */
  assign n1262_o = opc_opcode_q == 8'b01011010;
  /* decoder_pack-p.vhd:138:36  */
  assign n1263_o = n1260_o | n1262_o;
  /* decoder_pack-p.vhd:138:49  */
  assign n1265_o = opc_opcode_q == 8'b01011011;
  /* decoder_pack-p.vhd:138:49  */
  assign n1266_o = n1263_o | n1265_o;
  /* decoder_pack-p.vhd:138:62  */
  assign n1268_o = opc_opcode_q == 8'b01011100;
  /* decoder_pack-p.vhd:138:62  */
  assign n1269_o = n1266_o | n1268_o;
  /* decoder_pack-p.vhd:139:23  */
  assign n1271_o = opc_opcode_q == 8'b01011101;
  /* decoder_pack-p.vhd:139:23  */
  assign n1272_o = n1269_o | n1271_o;
  /* decoder_pack-p.vhd:139:36  */
  assign n1274_o = opc_opcode_q == 8'b01011110;
  /* decoder_pack-p.vhd:139:36  */
  assign n1275_o = n1272_o | n1274_o;
  /* decoder_pack-p.vhd:139:49  */
  assign n1277_o = opc_opcode_q == 8'b01011111;
  /* decoder_pack-p.vhd:139:49  */
  assign n1278_o = n1275_o | n1277_o;
  /* decoder_pack-p.vhd:139:62  */
  assign n1280_o = opc_opcode_q == 8'b01010000;
  /* decoder_pack-p.vhd:139:62  */
  assign n1281_o = n1278_o | n1280_o;
  /* decoder_pack-p.vhd:140:23  */
  assign n1283_o = opc_opcode_q == 8'b01010001;
  /* decoder_pack-p.vhd:140:23  */
  assign n1284_o = n1281_o | n1283_o;
  /* decoder_pack-p.vhd:144:7  */
  assign n1286_o = opc_opcode_q == 8'b01010011;
  /* decoder_pack-p.vhd:149:7  */
  assign n1288_o = opc_opcode_q == 8'b00010100;
  /* decoder_pack-p.vhd:149:23  */
  assign n1290_o = opc_opcode_q == 8'b00110100;
  /* decoder_pack-p.vhd:149:23  */
  assign n1291_o = n1288_o | n1290_o;
  /* decoder_pack-p.vhd:149:36  */
  assign n1293_o = opc_opcode_q == 8'b01010100;
  /* decoder_pack-p.vhd:149:36  */
  assign n1294_o = n1291_o | n1293_o;
  /* decoder_pack-p.vhd:149:49  */
  assign n1296_o = opc_opcode_q == 8'b01110100;
  /* decoder_pack-p.vhd:149:49  */
  assign n1297_o = n1294_o | n1296_o;
  /* decoder_pack-p.vhd:149:62  */
  assign n1299_o = opc_opcode_q == 8'b10010100;
  /* decoder_pack-p.vhd:149:62  */
  assign n1300_o = n1297_o | n1299_o;
  /* decoder_pack-p.vhd:150:23  */
  assign n1302_o = opc_opcode_q == 8'b10110100;
  /* decoder_pack-p.vhd:150:23  */
  assign n1303_o = n1300_o | n1302_o;
  /* decoder_pack-p.vhd:150:36  */
  assign n1305_o = opc_opcode_q == 8'b11010100;
  /* decoder_pack-p.vhd:150:36  */
  assign n1306_o = n1303_o | n1305_o;
  /* decoder_pack-p.vhd:150:49  */
  assign n1308_o = opc_opcode_q == 8'b11110100;
  /* decoder_pack-p.vhd:150:49  */
  assign n1309_o = n1306_o | n1308_o;
  /* decoder_pack-p.vhd:155:7  */
  assign n1311_o = opc_opcode_q == 8'b00100111;
  /* decoder_pack-p.vhd:159:7  */
  assign n1313_o = opc_opcode_q == 8'b10010111;
  /* decoder_pack-p.vhd:163:7  */
  assign n1315_o = opc_opcode_q == 8'b10000101;
  /* decoder_pack-p.vhd:163:23  */
  assign n1317_o = opc_opcode_q == 8'b10100101;
  /* decoder_pack-p.vhd:163:23  */
  assign n1318_o = n1315_o | n1317_o;
  /* decoder_pack-p.vhd:168:7  */
  assign n1320_o = opc_opcode_q == 8'b00110111;
  /* decoder_pack-p.vhd:172:7  */
  assign n1322_o = opc_opcode_q == 8'b10100111;
  /* decoder_pack-p.vhd:176:7  */
  assign n1324_o = opc_opcode_q == 8'b10010101;
  /* decoder_pack-p.vhd:176:23  */
  assign n1326_o = opc_opcode_q == 8'b10110101;
  /* decoder_pack-p.vhd:176:23  */
  assign n1327_o = n1324_o | n1326_o;
  /* decoder_pack-p.vhd:181:7  */
  assign n1329_o = opc_opcode_q == 8'b01010111;
  /* decoder_pack-p.vhd:185:7  */
  assign n1331_o = opc_opcode_q == 8'b11001000;
  /* decoder_pack-p.vhd:185:23  */
  assign n1333_o = opc_opcode_q == 8'b11001001;
  /* decoder_pack-p.vhd:185:23  */
  assign n1334_o = n1331_o | n1333_o;
  /* decoder_pack-p.vhd:185:36  */
  assign n1336_o = opc_opcode_q == 8'b11001010;
  /* decoder_pack-p.vhd:185:36  */
  assign n1337_o = n1334_o | n1336_o;
  /* decoder_pack-p.vhd:185:49  */
  assign n1339_o = opc_opcode_q == 8'b11001011;
  /* decoder_pack-p.vhd:185:49  */
  assign n1340_o = n1337_o | n1339_o;
  /* decoder_pack-p.vhd:185:62  */
  assign n1342_o = opc_opcode_q == 8'b11001100;
  /* decoder_pack-p.vhd:185:62  */
  assign n1343_o = n1340_o | n1342_o;
  /* decoder_pack-p.vhd:186:23  */
  assign n1345_o = opc_opcode_q == 8'b11001101;
  /* decoder_pack-p.vhd:186:23  */
  assign n1346_o = n1343_o | n1345_o;
  /* decoder_pack-p.vhd:186:36  */
  assign n1348_o = opc_opcode_q == 8'b11001110;
  /* decoder_pack-p.vhd:186:36  */
  assign n1349_o = n1346_o | n1348_o;
  /* decoder_pack-p.vhd:186:49  */
  assign n1351_o = opc_opcode_q == 8'b11001111;
  /* decoder_pack-p.vhd:186:49  */
  assign n1352_o = n1349_o | n1351_o;
  /* decoder_pack-p.vhd:186:62  */
  assign n1354_o = opc_opcode_q == 8'b00000111;
  /* decoder_pack-p.vhd:186:62  */
  assign n1355_o = n1352_o | n1354_o;
  /* decoder_pack-p.vhd:191:7  */
  assign n1357_o = opc_opcode_q == 8'b00010101;
  /* decoder_pack-p.vhd:191:23  */
  assign n1359_o = opc_opcode_q == 8'b00000101;
  /* decoder_pack-p.vhd:191:23  */
  assign n1360_o = n1357_o | n1359_o;
  /* decoder_pack-p.vhd:196:7  */
  assign n1362_o = opc_opcode_q == 8'b00110101;
  /* decoder_pack-p.vhd:196:23  */
  assign n1364_o = opc_opcode_q == 8'b00100101;
  /* decoder_pack-p.vhd:196:23  */
  assign n1365_o = n1362_o | n1364_o;
  /* decoder_pack-p.vhd:201:7  */
  assign n1367_o = opc_opcode_q == 8'b11101000;
  /* decoder_pack-p.vhd:201:23  */
  assign n1369_o = opc_opcode_q == 8'b11101001;
  /* decoder_pack-p.vhd:201:23  */
  assign n1370_o = n1367_o | n1369_o;
  /* decoder_pack-p.vhd:201:36  */
  assign n1372_o = opc_opcode_q == 8'b11101010;
  /* decoder_pack-p.vhd:201:36  */
  assign n1373_o = n1370_o | n1372_o;
  /* decoder_pack-p.vhd:201:49  */
  assign n1375_o = opc_opcode_q == 8'b11101011;
  /* decoder_pack-p.vhd:201:49  */
  assign n1376_o = n1373_o | n1375_o;
  /* decoder_pack-p.vhd:201:62  */
  assign n1378_o = opc_opcode_q == 8'b11101100;
  /* decoder_pack-p.vhd:201:62  */
  assign n1379_o = n1376_o | n1378_o;
  /* decoder_pack-p.vhd:202:23  */
  assign n1381_o = opc_opcode_q == 8'b11101101;
  /* decoder_pack-p.vhd:202:23  */
  assign n1382_o = n1379_o | n1381_o;
  /* decoder_pack-p.vhd:202:36  */
  assign n1384_o = opc_opcode_q == 8'b11101110;
  /* decoder_pack-p.vhd:202:36  */
  assign n1385_o = n1382_o | n1384_o;
  /* decoder_pack-p.vhd:202:49  */
  assign n1387_o = opc_opcode_q == 8'b11101111;
  /* decoder_pack-p.vhd:202:49  */
  assign n1388_o = n1385_o | n1387_o;
  /* decoder_pack-p.vhd:207:7  */
  assign n1390_o = opc_opcode_q == 8'b00001001;
  /* decoder_pack-p.vhd:207:23  */
  assign n1392_o = opc_opcode_q == 8'b00001010;
  /* decoder_pack-p.vhd:207:23  */
  assign n1393_o = n1390_o | n1392_o;
  /* decoder_pack-p.vhd:212:7  */
  assign n1395_o = opc_opcode_q == 8'b00010111;
  /* decoder_pack-p.vhd:212:23  */
  assign n1397_o = opc_opcode_q == 8'b00011000;
  /* decoder_pack-p.vhd:212:23  */
  assign n1398_o = n1395_o | n1397_o;
  /* decoder_pack-p.vhd:213:23  */
  assign n1400_o = opc_opcode_q == 8'b00011001;
  /* decoder_pack-p.vhd:213:23  */
  assign n1401_o = n1398_o | n1400_o;
  /* decoder_pack-p.vhd:213:36  */
  assign n1403_o = opc_opcode_q == 8'b00011010;
  /* decoder_pack-p.vhd:213:36  */
  assign n1404_o = n1401_o | n1403_o;
  /* decoder_pack-p.vhd:213:49  */
  assign n1406_o = opc_opcode_q == 8'b00011011;
  /* decoder_pack-p.vhd:213:49  */
  assign n1407_o = n1404_o | n1406_o;
  /* decoder_pack-p.vhd:213:62  */
  assign n1409_o = opc_opcode_q == 8'b00011100;
  /* decoder_pack-p.vhd:213:62  */
  assign n1410_o = n1407_o | n1409_o;
  /* decoder_pack-p.vhd:214:23  */
  assign n1412_o = opc_opcode_q == 8'b00011101;
  /* decoder_pack-p.vhd:214:23  */
  assign n1413_o = n1410_o | n1412_o;
  /* decoder_pack-p.vhd:214:36  */
  assign n1415_o = opc_opcode_q == 8'b00011110;
  /* decoder_pack-p.vhd:214:36  */
  assign n1416_o = n1413_o | n1415_o;
  /* decoder_pack-p.vhd:214:49  */
  assign n1418_o = opc_opcode_q == 8'b00011111;
  /* decoder_pack-p.vhd:214:49  */
  assign n1419_o = n1416_o | n1418_o;
  /* decoder_pack-p.vhd:214:62  */
  assign n1421_o = opc_opcode_q == 8'b00010000;
  /* decoder_pack-p.vhd:214:62  */
  assign n1422_o = n1419_o | n1421_o;
  /* decoder_pack-p.vhd:215:23  */
  assign n1424_o = opc_opcode_q == 8'b00010001;
  /* decoder_pack-p.vhd:215:23  */
  assign n1425_o = n1422_o | n1424_o;
  /* decoder_pack-p.vhd:219:7  */
  assign n1427_o = opc_opcode_q == 8'b00010010;
  /* decoder_pack-p.vhd:219:23  */
  assign n1429_o = opc_opcode_q == 8'b00110010;
  /* decoder_pack-p.vhd:219:23  */
  assign n1430_o = n1427_o | n1429_o;
  /* decoder_pack-p.vhd:219:36  */
  assign n1432_o = opc_opcode_q == 8'b01010010;
  /* decoder_pack-p.vhd:219:36  */
  assign n1433_o = n1430_o | n1432_o;
  /* decoder_pack-p.vhd:219:49  */
  assign n1435_o = opc_opcode_q == 8'b01110010;
  /* decoder_pack-p.vhd:219:49  */
  assign n1436_o = n1433_o | n1435_o;
  /* decoder_pack-p.vhd:219:62  */
  assign n1438_o = opc_opcode_q == 8'b10010010;
  /* decoder_pack-p.vhd:219:62  */
  assign n1439_o = n1436_o | n1438_o;
  /* decoder_pack-p.vhd:220:23  */
  assign n1441_o = opc_opcode_q == 8'b10110010;
  /* decoder_pack-p.vhd:220:23  */
  assign n1442_o = n1439_o | n1441_o;
  /* decoder_pack-p.vhd:220:36  */
  assign n1444_o = opc_opcode_q == 8'b11010010;
  /* decoder_pack-p.vhd:220:36  */
  assign n1445_o = n1442_o | n1444_o;
  /* decoder_pack-p.vhd:220:49  */
  assign n1447_o = opc_opcode_q == 8'b11110010;
  /* decoder_pack-p.vhd:220:49  */
  assign n1448_o = n1445_o | n1447_o;
  /* decoder_pack-p.vhd:225:7  */
  assign n1450_o = opc_opcode_q == 8'b11110110;
  /* decoder_pack-p.vhd:225:23  */
  assign n1452_o = opc_opcode_q == 8'b11100110;
  /* decoder_pack-p.vhd:225:23  */
  assign n1453_o = n1450_o | n1452_o;
  /* decoder_pack-p.vhd:231:7  */
  assign n1455_o = opc_opcode_q == 8'b10110110;
  /* decoder_pack-p.vhd:231:23  */
  assign n1457_o = opc_opcode_q == 8'b01110110;
  /* decoder_pack-p.vhd:231:23  */
  assign n1458_o = n1455_o | n1457_o;
  /* decoder_pack-p.vhd:237:7  */
  assign n1460_o = opc_opcode_q == 8'b00000100;
  /* decoder_pack-p.vhd:237:23  */
  assign n1462_o = opc_opcode_q == 8'b00100100;
  /* decoder_pack-p.vhd:237:23  */
  assign n1463_o = n1460_o | n1462_o;
  /* decoder_pack-p.vhd:237:36  */
  assign n1465_o = opc_opcode_q == 8'b01000100;
  /* decoder_pack-p.vhd:237:36  */
  assign n1466_o = n1463_o | n1465_o;
  /* decoder_pack-p.vhd:237:49  */
  assign n1468_o = opc_opcode_q == 8'b01100100;
  /* decoder_pack-p.vhd:237:49  */
  assign n1469_o = n1466_o | n1468_o;
  /* decoder_pack-p.vhd:237:62  */
  assign n1471_o = opc_opcode_q == 8'b10000100;
  /* decoder_pack-p.vhd:237:62  */
  assign n1472_o = n1469_o | n1471_o;
  /* decoder_pack-p.vhd:238:23  */
  assign n1474_o = opc_opcode_q == 8'b10100100;
  /* decoder_pack-p.vhd:238:23  */
  assign n1475_o = n1472_o | n1474_o;
  /* decoder_pack-p.vhd:238:36  */
  assign n1477_o = opc_opcode_q == 8'b11000100;
  /* decoder_pack-p.vhd:238:36  */
  assign n1478_o = n1475_o | n1477_o;
  /* decoder_pack-p.vhd:238:49  */
  assign n1480_o = opc_opcode_q == 8'b11100100;
  /* decoder_pack-p.vhd:238:49  */
  assign n1481_o = n1478_o | n1480_o;
  /* decoder_pack-p.vhd:243:7  */
  assign n1483_o = opc_opcode_q == 8'b10110011;
  /* decoder_pack-p.vhd:248:7  */
  assign n1485_o = opc_opcode_q == 8'b00100110;
  /* decoder_pack-p.vhd:248:23  */
  assign n1487_o = opc_opcode_q == 8'b01000110;
  /* decoder_pack-p.vhd:248:23  */
  assign n1488_o = n1485_o | n1487_o;
  /* decoder_pack-p.vhd:249:23  */
  assign n1490_o = opc_opcode_q == 8'b00110110;
  /* decoder_pack-p.vhd:249:23  */
  assign n1491_o = n1488_o | n1490_o;
  /* decoder_pack-p.vhd:250:23  */
  assign n1493_o = opc_opcode_q == 8'b01010110;
  /* decoder_pack-p.vhd:250:23  */
  assign n1494_o = n1491_o | n1493_o;
  /* decoder_pack-p.vhd:256:7  */
  assign n1496_o = opc_opcode_q == 8'b00010110;
  /* decoder_pack-p.vhd:261:7  */
  assign n1498_o = opc_opcode_q == 8'b10010110;
  /* decoder_pack-p.vhd:261:23  */
  assign n1500_o = opc_opcode_q == 8'b11000110;
  /* decoder_pack-p.vhd:261:23  */
  assign n1501_o = n1498_o | n1500_o;
  /* decoder_pack-p.vhd:267:7  */
  assign n1503_o = opc_opcode_q == 8'b00100011;
  /* decoder_pack-p.vhd:272:7  */
  assign n1505_o = opc_opcode_q == 8'b11000111;
  /* decoder_pack-p.vhd:276:7  */
  assign n1507_o = opc_opcode_q == 8'b11111000;
  /* decoder_pack-p.vhd:276:23  */
  assign n1509_o = opc_opcode_q == 8'b11111001;
  /* decoder_pack-p.vhd:276:23  */
  assign n1510_o = n1507_o | n1509_o;
  /* decoder_pack-p.vhd:276:36  */
  assign n1512_o = opc_opcode_q == 8'b11111010;
  /* decoder_pack-p.vhd:276:36  */
  assign n1513_o = n1510_o | n1512_o;
  /* decoder_pack-p.vhd:276:49  */
  assign n1515_o = opc_opcode_q == 8'b11111011;
  /* decoder_pack-p.vhd:276:49  */
  assign n1516_o = n1513_o | n1515_o;
  /* decoder_pack-p.vhd:276:62  */
  assign n1518_o = opc_opcode_q == 8'b11111100;
  /* decoder_pack-p.vhd:276:62  */
  assign n1519_o = n1516_o | n1518_o;
  /* decoder_pack-p.vhd:277:23  */
  assign n1521_o = opc_opcode_q == 8'b11111101;
  /* decoder_pack-p.vhd:277:23  */
  assign n1522_o = n1519_o | n1521_o;
  /* decoder_pack-p.vhd:277:36  */
  assign n1524_o = opc_opcode_q == 8'b11111110;
  /* decoder_pack-p.vhd:277:36  */
  assign n1525_o = n1522_o | n1524_o;
  /* decoder_pack-p.vhd:277:49  */
  assign n1527_o = opc_opcode_q == 8'b11111111;
  /* decoder_pack-p.vhd:277:49  */
  assign n1528_o = n1525_o | n1527_o;
  /* decoder_pack-p.vhd:277:62  */
  assign n1530_o = opc_opcode_q == 8'b11110000;
  /* decoder_pack-p.vhd:277:62  */
  assign n1531_o = n1528_o | n1530_o;
  /* decoder_pack-p.vhd:278:23  */
  assign n1533_o = opc_opcode_q == 8'b11110001;
  /* decoder_pack-p.vhd:278:23  */
  assign n1534_o = n1531_o | n1533_o;
  /* decoder_pack-p.vhd:282:7  */
  assign n1536_o = opc_opcode_q == 8'b11010111;
  /* decoder_pack-p.vhd:286:7  */
  assign n1538_o = opc_opcode_q == 8'b10101000;
  /* decoder_pack-p.vhd:286:23  */
  assign n1540_o = opc_opcode_q == 8'b10101001;
  /* decoder_pack-p.vhd:286:23  */
  assign n1541_o = n1538_o | n1540_o;
  /* decoder_pack-p.vhd:286:36  */
  assign n1543_o = opc_opcode_q == 8'b10101010;
  /* decoder_pack-p.vhd:286:36  */
  assign n1544_o = n1541_o | n1543_o;
  /* decoder_pack-p.vhd:286:49  */
  assign n1546_o = opc_opcode_q == 8'b10101011;
  /* decoder_pack-p.vhd:286:49  */
  assign n1547_o = n1544_o | n1546_o;
  /* decoder_pack-p.vhd:286:62  */
  assign n1549_o = opc_opcode_q == 8'b10101100;
  /* decoder_pack-p.vhd:286:62  */
  assign n1550_o = n1547_o | n1549_o;
  /* decoder_pack-p.vhd:287:23  */
  assign n1552_o = opc_opcode_q == 8'b10101101;
  /* decoder_pack-p.vhd:287:23  */
  assign n1553_o = n1550_o | n1552_o;
  /* decoder_pack-p.vhd:287:36  */
  assign n1555_o = opc_opcode_q == 8'b10101110;
  /* decoder_pack-p.vhd:287:36  */
  assign n1556_o = n1553_o | n1555_o;
  /* decoder_pack-p.vhd:287:49  */
  assign n1558_o = opc_opcode_q == 8'b10101111;
  /* decoder_pack-p.vhd:287:49  */
  assign n1559_o = n1556_o | n1558_o;
  /* decoder_pack-p.vhd:287:62  */
  assign n1561_o = opc_opcode_q == 8'b10100000;
  /* decoder_pack-p.vhd:287:62  */
  assign n1562_o = n1559_o | n1561_o;
  /* decoder_pack-p.vhd:288:23  */
  assign n1564_o = opc_opcode_q == 8'b10100001;
  /* decoder_pack-p.vhd:288:23  */
  assign n1565_o = n1562_o | n1564_o;
  /* decoder_pack-p.vhd:292:7  */
  assign n1567_o = opc_opcode_q == 8'b10111000;
  /* decoder_pack-p.vhd:292:23  */
  assign n1569_o = opc_opcode_q == 8'b10111001;
  /* decoder_pack-p.vhd:292:23  */
  assign n1570_o = n1567_o | n1569_o;
  /* decoder_pack-p.vhd:292:36  */
  assign n1572_o = opc_opcode_q == 8'b10111010;
  /* decoder_pack-p.vhd:292:36  */
  assign n1573_o = n1570_o | n1572_o;
  /* decoder_pack-p.vhd:292:49  */
  assign n1575_o = opc_opcode_q == 8'b10111011;
  /* decoder_pack-p.vhd:292:49  */
  assign n1576_o = n1573_o | n1575_o;
  /* decoder_pack-p.vhd:292:62  */
  assign n1578_o = opc_opcode_q == 8'b10111100;
  /* decoder_pack-p.vhd:292:62  */
  assign n1579_o = n1576_o | n1578_o;
  /* decoder_pack-p.vhd:293:23  */
  assign n1581_o = opc_opcode_q == 8'b10111101;
  /* decoder_pack-p.vhd:293:23  */
  assign n1582_o = n1579_o | n1581_o;
  /* decoder_pack-p.vhd:293:36  */
  assign n1584_o = opc_opcode_q == 8'b10111110;
  /* decoder_pack-p.vhd:293:36  */
  assign n1585_o = n1582_o | n1584_o;
  /* decoder_pack-p.vhd:293:49  */
  assign n1587_o = opc_opcode_q == 8'b10111111;
  /* decoder_pack-p.vhd:293:49  */
  assign n1588_o = n1585_o | n1587_o;
  /* decoder_pack-p.vhd:293:62  */
  assign n1590_o = opc_opcode_q == 8'b10110000;
  /* decoder_pack-p.vhd:293:62  */
  assign n1591_o = n1588_o | n1590_o;
  /* decoder_pack-p.vhd:294:23  */
  assign n1593_o = opc_opcode_q == 8'b10110001;
  /* decoder_pack-p.vhd:294:23  */
  assign n1594_o = n1591_o | n1593_o;
  /* decoder_pack-p.vhd:299:7  */
  assign n1596_o = opc_opcode_q == 8'b01100010;
  /* decoder_pack-p.vhd:299:23  */
  assign n1598_o = opc_opcode_q == 8'b01000010;
  /* decoder_pack-p.vhd:299:23  */
  assign n1599_o = n1596_o | n1598_o;
  /* decoder_pack-p.vhd:304:7  */
  assign n1601_o = opc_opcode_q == 8'b00001100;
  /* decoder_pack-p.vhd:304:23  */
  assign n1603_o = opc_opcode_q == 8'b00001101;
  /* decoder_pack-p.vhd:304:23  */
  assign n1604_o = n1601_o | n1603_o;
  /* decoder_pack-p.vhd:304:36  */
  assign n1606_o = opc_opcode_q == 8'b00001110;
  /* decoder_pack-p.vhd:304:36  */
  assign n1607_o = n1604_o | n1606_o;
  /* decoder_pack-p.vhd:304:49  */
  assign n1609_o = opc_opcode_q == 8'b00001111;
  /* decoder_pack-p.vhd:304:49  */
  assign n1610_o = n1607_o | n1609_o;
  /* decoder_pack-p.vhd:309:7  */
  assign n1612_o = opc_opcode_q == 8'b10100011;
  /* decoder_pack-p.vhd:309:23  */
  assign n1614_o = opc_opcode_q == 8'b11100011;
  /* decoder_pack-p.vhd:309:23  */
  assign n1615_o = n1612_o | n1614_o;
  /* decoder_pack-p.vhd:315:7  */
  assign n1617_o = opc_opcode_q == 8'b00000000;
  /* decoder_pack-p.vhd:319:7  */
  assign n1619_o = opc_opcode_q == 8'b01001000;
  /* decoder_pack-p.vhd:319:23  */
  assign n1621_o = opc_opcode_q == 8'b01001001;
  /* decoder_pack-p.vhd:319:23  */
  assign n1622_o = n1619_o | n1621_o;
  /* decoder_pack-p.vhd:319:36  */
  assign n1624_o = opc_opcode_q == 8'b01001010;
  /* decoder_pack-p.vhd:319:36  */
  assign n1625_o = n1622_o | n1624_o;
  /* decoder_pack-p.vhd:319:49  */
  assign n1627_o = opc_opcode_q == 8'b01001011;
  /* decoder_pack-p.vhd:319:49  */
  assign n1628_o = n1625_o | n1627_o;
  /* decoder_pack-p.vhd:319:62  */
  assign n1630_o = opc_opcode_q == 8'b01001100;
  /* decoder_pack-p.vhd:319:62  */
  assign n1631_o = n1628_o | n1630_o;
  /* decoder_pack-p.vhd:320:23  */
  assign n1633_o = opc_opcode_q == 8'b01001101;
  /* decoder_pack-p.vhd:320:23  */
  assign n1634_o = n1631_o | n1633_o;
  /* decoder_pack-p.vhd:320:36  */
  assign n1636_o = opc_opcode_q == 8'b01001110;
  /* decoder_pack-p.vhd:320:36  */
  assign n1637_o = n1634_o | n1636_o;
  /* decoder_pack-p.vhd:320:49  */
  assign n1639_o = opc_opcode_q == 8'b01001111;
  /* decoder_pack-p.vhd:320:49  */
  assign n1640_o = n1637_o | n1639_o;
  /* decoder_pack-p.vhd:320:62  */
  assign n1642_o = opc_opcode_q == 8'b01000000;
  /* decoder_pack-p.vhd:320:62  */
  assign n1643_o = n1640_o | n1642_o;
  /* decoder_pack-p.vhd:321:23  */
  assign n1645_o = opc_opcode_q == 8'b01000001;
  /* decoder_pack-p.vhd:321:23  */
  assign n1646_o = n1643_o | n1645_o;
  /* decoder_pack-p.vhd:325:7  */
  assign n1648_o = opc_opcode_q == 8'b01000011;
  /* decoder_pack-p.vhd:330:7  */
  assign n1650_o = opc_opcode_q == 8'b00111100;
  /* decoder_pack-p.vhd:330:23  */
  assign n1652_o = opc_opcode_q == 8'b00111101;
  /* decoder_pack-p.vhd:330:23  */
  assign n1653_o = n1650_o | n1652_o;
  /* decoder_pack-p.vhd:330:36  */
  assign n1655_o = opc_opcode_q == 8'b00111110;
  /* decoder_pack-p.vhd:330:36  */
  assign n1656_o = n1653_o | n1655_o;
  /* decoder_pack-p.vhd:330:49  */
  assign n1658_o = opc_opcode_q == 8'b00111111;
  /* decoder_pack-p.vhd:330:49  */
  assign n1659_o = n1656_o | n1658_o;
  /* decoder_pack-p.vhd:330:62  */
  assign n1661_o = opc_opcode_q == 8'b10011100;
  /* decoder_pack-p.vhd:330:62  */
  assign n1662_o = n1659_o | n1661_o;
  /* decoder_pack-p.vhd:331:23  */
  assign n1664_o = opc_opcode_q == 8'b10011101;
  /* decoder_pack-p.vhd:331:23  */
  assign n1665_o = n1662_o | n1664_o;
  /* decoder_pack-p.vhd:331:36  */
  assign n1667_o = opc_opcode_q == 8'b10011110;
  /* decoder_pack-p.vhd:331:36  */
  assign n1668_o = n1665_o | n1667_o;
  /* decoder_pack-p.vhd:331:49  */
  assign n1670_o = opc_opcode_q == 8'b10011111;
  /* decoder_pack-p.vhd:331:49  */
  assign n1671_o = n1668_o | n1670_o;
  /* decoder_pack-p.vhd:331:62  */
  assign n1673_o = opc_opcode_q == 8'b10001100;
  /* decoder_pack-p.vhd:331:62  */
  assign n1674_o = n1671_o | n1673_o;
  /* decoder_pack-p.vhd:332:23  */
  assign n1676_o = opc_opcode_q == 8'b10001101;
  /* decoder_pack-p.vhd:332:23  */
  assign n1677_o = n1674_o | n1676_o;
  /* decoder_pack-p.vhd:332:36  */
  assign n1679_o = opc_opcode_q == 8'b10001110;
  /* decoder_pack-p.vhd:332:36  */
  assign n1680_o = n1677_o | n1679_o;
  /* decoder_pack-p.vhd:332:49  */
  assign n1682_o = opc_opcode_q == 8'b10001111;
  /* decoder_pack-p.vhd:332:49  */
  assign n1683_o = n1680_o | n1682_o;
  /* decoder_pack-p.vhd:337:7  */
  assign n1685_o = opc_opcode_q == 8'b10000011;
  /* decoder_pack-p.vhd:337:23  */
  assign n1687_o = opc_opcode_q == 8'b10010011;
  /* decoder_pack-p.vhd:337:23  */
  assign n1688_o = n1685_o | n1687_o;
  /* decoder_pack-p.vhd:343:7  */
  assign n1690_o = opc_opcode_q == 8'b11100111;
  /* decoder_pack-p.vhd:343:23  */
  assign n1692_o = opc_opcode_q == 8'b11110111;
  /* decoder_pack-p.vhd:343:23  */
  assign n1693_o = n1690_o | n1692_o;
  /* decoder_pack-p.vhd:348:7  */
  assign n1695_o = opc_opcode_q == 8'b01110111;
  /* decoder_pack-p.vhd:348:23  */
  assign n1697_o = opc_opcode_q == 8'b01100111;
  /* decoder_pack-p.vhd:348:23  */
  assign n1698_o = n1695_o | n1697_o;
  /* decoder_pack-p.vhd:353:7  */
  assign n1700_o = opc_opcode_q == 8'b11000101;
  /* decoder_pack-p.vhd:353:23  */
  assign n1702_o = opc_opcode_q == 8'b11010101;
  /* decoder_pack-p.vhd:353:23  */
  assign n1703_o = n1700_o | n1702_o;
  /* decoder_pack-p.vhd:358:7  */
  assign n1705_o = opc_opcode_q == 8'b01100101;
  /* decoder_pack-p.vhd:362:7  */
  assign n1707_o = opc_opcode_q == 8'b01000101;
  /* decoder_pack-p.vhd:362:23  */
  assign n1709_o = opc_opcode_q == 8'b01010101;
  /* decoder_pack-p.vhd:362:23  */
  assign n1710_o = n1707_o | n1709_o;
  /* decoder_pack-p.vhd:367:7  */
  assign n1712_o = opc_opcode_q == 8'b01000111;
  /* decoder_pack-p.vhd:371:7  */
  assign n1714_o = opc_opcode_q == 8'b00101000;
  /* decoder_pack-p.vhd:371:23  */
  assign n1716_o = opc_opcode_q == 8'b00101001;
  /* decoder_pack-p.vhd:371:23  */
  assign n1717_o = n1714_o | n1716_o;
  /* decoder_pack-p.vhd:371:36  */
  assign n1719_o = opc_opcode_q == 8'b00101010;
  /* decoder_pack-p.vhd:371:36  */
  assign n1720_o = n1717_o | n1719_o;
  /* decoder_pack-p.vhd:371:49  */
  assign n1722_o = opc_opcode_q == 8'b00101011;
  /* decoder_pack-p.vhd:371:49  */
  assign n1723_o = n1720_o | n1722_o;
  /* decoder_pack-p.vhd:371:62  */
  assign n1725_o = opc_opcode_q == 8'b00101100;
  /* decoder_pack-p.vhd:371:62  */
  assign n1726_o = n1723_o | n1725_o;
  /* decoder_pack-p.vhd:372:23  */
  assign n1728_o = opc_opcode_q == 8'b00101101;
  /* decoder_pack-p.vhd:372:23  */
  assign n1729_o = n1726_o | n1728_o;
  /* decoder_pack-p.vhd:372:36  */
  assign n1731_o = opc_opcode_q == 8'b00101110;
  /* decoder_pack-p.vhd:372:36  */
  assign n1732_o = n1729_o | n1731_o;
  /* decoder_pack-p.vhd:372:49  */
  assign n1734_o = opc_opcode_q == 8'b00101111;
  /* decoder_pack-p.vhd:372:49  */
  assign n1735_o = n1732_o | n1734_o;
  /* decoder_pack-p.vhd:372:62  */
  assign n1737_o = opc_opcode_q == 8'b00100000;
  /* decoder_pack-p.vhd:372:62  */
  assign n1738_o = n1735_o | n1737_o;
  /* decoder_pack-p.vhd:373:23  */
  assign n1740_o = opc_opcode_q == 8'b00100001;
  /* decoder_pack-p.vhd:373:23  */
  assign n1741_o = n1738_o | n1740_o;
  /* decoder_pack-p.vhd:373:36  */
  assign n1743_o = opc_opcode_q == 8'b00110000;
  /* decoder_pack-p.vhd:373:36  */
  assign n1744_o = n1741_o | n1743_o;
  /* decoder_pack-p.vhd:374:23  */
  assign n1746_o = opc_opcode_q == 8'b00110001;
  /* decoder_pack-p.vhd:374:23  */
  assign n1747_o = n1744_o | n1746_o;
  /* decoder_pack-p.vhd:378:7  */
  assign n1749_o = opc_opcode_q == 8'b11011000;
  /* decoder_pack-p.vhd:378:23  */
  assign n1751_o = opc_opcode_q == 8'b11011001;
  /* decoder_pack-p.vhd:378:23  */
  assign n1752_o = n1749_o | n1751_o;
  /* decoder_pack-p.vhd:378:36  */
  assign n1754_o = opc_opcode_q == 8'b11011010;
  /* decoder_pack-p.vhd:378:36  */
  assign n1755_o = n1752_o | n1754_o;
  /* decoder_pack-p.vhd:378:49  */
  assign n1757_o = opc_opcode_q == 8'b11011011;
  /* decoder_pack-p.vhd:378:49  */
  assign n1758_o = n1755_o | n1757_o;
  /* decoder_pack-p.vhd:378:62  */
  assign n1760_o = opc_opcode_q == 8'b11011100;
  /* decoder_pack-p.vhd:378:62  */
  assign n1761_o = n1758_o | n1760_o;
  /* decoder_pack-p.vhd:379:23  */
  assign n1763_o = opc_opcode_q == 8'b11011101;
  /* decoder_pack-p.vhd:379:23  */
  assign n1764_o = n1761_o | n1763_o;
  /* decoder_pack-p.vhd:379:36  */
  assign n1766_o = opc_opcode_q == 8'b11011110;
  /* decoder_pack-p.vhd:379:36  */
  assign n1767_o = n1764_o | n1766_o;
  /* decoder_pack-p.vhd:379:49  */
  assign n1769_o = opc_opcode_q == 8'b11011111;
  /* decoder_pack-p.vhd:379:49  */
  assign n1770_o = n1767_o | n1769_o;
  /* decoder_pack-p.vhd:379:62  */
  assign n1772_o = opc_opcode_q == 8'b11010000;
  /* decoder_pack-p.vhd:379:62  */
  assign n1773_o = n1770_o | n1772_o;
  /* decoder_pack-p.vhd:380:23  */
  assign n1775_o = opc_opcode_q == 8'b11010001;
  /* decoder_pack-p.vhd:380:23  */
  assign n1776_o = n1773_o | n1775_o;
  /* decoder_pack-p.vhd:384:7  */
  assign n1778_o = opc_opcode_q == 8'b11010011;
  assign n1779_o = {n1778_o, n1776_o, n1747_o, n1712_o, n1710_o, n1705_o, n1703_o, n1698_o, n1693_o, n1688_o, n1683_o, n1648_o, n1646_o, n1617_o, n1615_o, n1610_o, n1599_o, n1594_o, n1565_o, n1536_o, n1534_o, n1505_o, n1503_o, n1501_o, n1496_o, n1494_o, n1483_o, n1481_o, n1458_o, n1453_o, n1448_o, n1425_o, n1393_o, n1388_o, n1365_o, n1360_o, n1355_o, n1329_o, n1327_o, n1322_o, n1320_o, n1318_o, n1313_o, n1311_o, n1309_o, n1286_o, n1284_o, n1255_o, n1250_o};
  /* decoder_pack-p.vhd:121:5  */
  always @*
    case (n1779_o)
      49'b1000000000000000000000000000000000000000000000000: n1830_o = 6'b111001;
      49'b0100000000000000000000000000000000000000000000000: n1830_o = 6'b111000;
      49'b0010000000000000000000000000000000000000000000000: n1830_o = 6'b110111;
      49'b0001000000000000000000000000000000000000000000000: n1830_o = 6'b110110;
      49'b0000100000000000000000000000000000000000000000000: n1830_o = 6'b110101;
      49'b0000010000000000000000000000000000000000000000000: n1830_o = 6'b110100;
      49'b0000001000000000000000000000000000000000000000000: n1830_o = 6'b110011;
      49'b0000000100000000000000000000000000000000000000000: n1830_o = 6'b110001;
      49'b0000000010000000000000000000000000000000000000000: n1830_o = 6'b110000;
      49'b0000000001000000000000000000000000000000000000000: n1830_o = 6'b101111;
      49'b0000000000100000000000000000000000000000000000000: n1830_o = 6'b101101;
      49'b0000000000010000000000000000000000000000000000000: n1830_o = 6'b101011;
      49'b0000000000001000000000000000000000000000000000000: n1830_o = 6'b101010;
      49'b0000000000000100000000000000000000000000000000000: n1830_o = 6'b101001;
      49'b0000000000000010000000000000000000000000000000000: n1830_o = 6'b100111;
      49'b0000000000000001000000000000000000000000000000000: n1830_o = 6'b100110;
      49'b0000000000000000100000000000000000000000000000000: n1830_o = 6'b100101;
      49'b0000000000000000010000000000000000000000000000000: n1830_o = 6'b100100;
      49'b0000000000000000001000000000000000000000000000000: n1830_o = 6'b100011;
      49'b0000000000000000000100000000000000000000000000000: n1830_o = 6'b100010;
      49'b0000000000000000000010000000000000000000000000000: n1830_o = 6'b100001;
      49'b0000000000000000000001000000000000000000000000000: n1830_o = 6'b100000;
      49'b0000000000000000000000100000000000000000000000000: n1830_o = 6'b011111;
      49'b0000000000000000000000010000000000000000000000000: n1830_o = 6'b011110;
      49'b0000000000000000000000001000000000000000000000000: n1830_o = 6'b011101;
      49'b0000000000000000000000000100000000000000000000000: n1830_o = 6'b011100;
      49'b0000000000000000000000000010000000000000000000000: n1830_o = 6'b011010;
      49'b0000000000000000000000000001000000000000000000000: n1830_o = 6'b011001;
      49'b0000000000000000000000000000100000000000000000000: n1830_o = 6'b011000;
      49'b0000000000000000000000000000010000000000000000000: n1830_o = 6'b010111;
      49'b0000000000000000000000000000001000000000000000000: n1830_o = 6'b010110;
      49'b0000000000000000000000000000000100000000000000000: n1830_o = 6'b010100;
      49'b0000000000000000000000000000000010000000000000000: n1830_o = 6'b010011;
      49'b0000000000000000000000000000000001000000000000000: n1830_o = 6'b010001;
      49'b0000000000000000000000000000000000100000000000000: n1830_o = 6'b010000;
      49'b0000000000000000000000000000000000010000000000000: n1830_o = 6'b001111;
      49'b0000000000000000000000000000000000001000000000000: n1830_o = 6'b001110;
      49'b0000000000000000000000000000000000000100000000000: n1830_o = 6'b001101;
      49'b0000000000000000000000000000000000000010000000000: n1830_o = 6'b001100;
      49'b0000000000000000000000000000000000000001000000000: n1830_o = 6'b001011;
      49'b0000000000000000000000000000000000000000100000000: n1830_o = 6'b001010;
      49'b0000000000000000000000000000000000000000010000000: n1830_o = 6'b001001;
      49'b0000000000000000000000000000000000000000001000000: n1830_o = 6'b001000;
      49'b0000000000000000000000000000000000000000000100000: n1830_o = 6'b000111;
      49'b0000000000000000000000000000000000000000000010000: n1830_o = 6'b000110;
      49'b0000000000000000000000000000000000000000000001000: n1830_o = 6'b000100;
      49'b0000000000000000000000000000000000000000000000100: n1830_o = 6'b000011;
      49'b0000000000000000000000000000000000000000000000010: n1830_o = 6'b000010;
      49'b0000000000000000000000000000000000000000000000001: n1830_o = 6'b000001;
      default: n1830_o = 6'b101001;
    endcase
  /* decoder_pack-p.vhd:121:5  */
  always @*
    case (n1779_o)
      49'b1000000000000000000000000000000000000000000000000: n1854_o = 1'b1;
      49'b0100000000000000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0010000000000000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0001000000000000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000100000000000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000010000000000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000001000000000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000100000000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000010000000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000001000000000000000000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000100000000000000000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000010000000000000000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000001000000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000000000100000000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000000000010000000000000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000001000000000000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000100000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000000000000010000000000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000001000000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000000000000000100000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000000000000000010000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000000000000000001000000000000000000000000000: n1854_o = 1'b0;
      49'b0000000000000000000000100000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000010000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000001000000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000100000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000010000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000001000000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000000100000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000000010000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000000001000000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000000000100000000000000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000010000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000000000001000000000000000: n1854_o = 1'b1;
      49'b0000000000000000000000000000000000100000000000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000010000000000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000001000000000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000100000000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000010000000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000001000000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000000100000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000000010000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000000001000000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000000000100000: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000000000010000: n1854_o = 1'b1;
      49'b0000000000000000000000000000000000000000000001000: n1854_o = 1'b1;
      49'b0000000000000000000000000000000000000000000000100: n1854_o = 1'b0;
      49'b0000000000000000000000000000000000000000000000010: n1854_o = 1'b1;
      49'b0000000000000000000000000000000000000000000000001: n1854_o = 1'b0;
      default: n1854_o = 1'b0;
    endcase
  assign n1858_o = {n1854_o, n1830_o};
  assign n1859_o = {n1180_o, n1171_o};
  /* decoder_pack-p.vhd:466:5  */
  assign n1860_o = n1183_o ? n1858_o : n1859_o;
  /* decoder.vhd:301:14  */
  assign n1863_o = ~res_i;
  /* decoder.vhd:313:40  */
  assign n1865_o = mnemonic_rec_s[5:0];
  /* decoder.vhd:310:9  */
  assign n1867_o = opc_inj_int_s ? 8'b00010100 : opc_opcode_q;
  /* decoder.vhd:310:9  */
  assign n1868_o = opc_inj_int_s ? mnemonic_q : n1865_o;
  /* decoder.vhd:308:9  */
  assign n1869_o = opc_read_bus_s ? data_i : n1867_o;
  /* decoder.vhd:308:9  */
  assign n1870_o = opc_read_bus_s ? mnemonic_q : n1868_o;
  /* decoder.vhd:322:39  */
  assign n1880_o = mnemonic_rec_s[6];
  /* decoder.vhd:324:24  */
  assign n1882_o = 1'b1 ? mnemonic_q : n1883_o;
  /* decoder.vhd:325:41  */
  assign n1883_o = mnemonic_rec_s[5:0];
  /* decoder.vhd:343:28  */
  assign int_b_n1884 = int_b_tf_o; // (signal)
  /* decoder.vhd:352:28  */
  assign int_b_n1886 = int_b_tim_int_o; // (signal)
  /* decoder.vhd:355:28  */
  assign int_b_n1887 = int_b_int_pending_o; // (signal)
  /* decoder.vhd:356:28  */
  assign int_b_n1888 = int_b_int_in_progress_o; // (signal)
  /* decoder.vhd:333:3  */
  t48_int int_b (
    .clk_i(clk_i),
    .res_i(res_i),
    .en_clk_i(en_clk_i),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_i),
    .clk_mstate_i(clk_mstate_i),
    .jtf_executed_i(jtf_executed_s),
    .tim_overflow_i(tim_overflow_i),
    .en_tcnti_i(en_tcnti_s),
    .dis_tcnti_i(dis_tcnti_s),
    .int_n_i(int_n_i),
    .ale_i(ale_i),
    .last_cycle_i(last_cycle_s),
    .en_i_i(en_i_s),
    .dis_i_i(dis_i_s),
    .retr_executed_i(retr_executed_s),
    .int_executed_i(int_executed_s),
    .tf_o(int_b_tf_o),
    .ext_int_o(),
    .tim_int_o(int_b_tim_int_o),
    .int_pending_o(int_b_int_pending_o),
    .int_in_progress_o(int_b_int_in_progress_o));
  /* decoder.vhd:359:19  */
  assign n1898_o = ~opc_multi_cycle_s;
  /* decoder.vhd:360:38  */
  assign n1899_o = clk_second_cycle_i & opc_multi_cycle_s;
  /* decoder.vhd:359:41  */
  assign n1900_o = n1898_o | n1899_o;
  /* decoder.vhd:393:26  */
  assign n1903_o = ~clk_second_cycle_i;
  /* decoder.vhd:394:46  */
  assign n1904_o = assert_psen_s & clk_second_cycle_i;
  /* decoder.vhd:393:49  */
  assign n1905_o = n1903_o | n1904_o;
  /* decoder.vhd:399:19  */
  assign n1906_o = ~ea_i;
  /* decoder.vhd:400:16  */
  assign n1907_o = ~int_pending_s;
  /* decoder.vhd:400:13  */
  assign n1910_o = n1907_o ? 1'b1 : 1'b0;
  /* decoder.vhd:405:16  */
  assign n1911_o = ~int_pending_s;
  /* decoder.vhd:405:13  */
  assign n1914_o = n1911_o ? 1'b1 : 1'b0;
  /* decoder.vhd:399:11  */
  assign n1916_o = n1906_o ? n1910_o : 1'b0;
  /* decoder.vhd:399:11  */
  assign n1919_o = n1906_o ? 1'b0 : 1'b1;
  /* decoder.vhd:399:11  */
  assign n1921_o = n1906_o ? 1'b0 : n1914_o;
  /* decoder.vhd:398:9  */
  assign n1923_o = n1905_o ? n1916_o : 1'b0;
  /* decoder.vhd:398:9  */
  assign n1925_o = n1905_o ? n1919_o : 1'b0;
  /* decoder.vhd:398:9  */
  assign n1927_o = n1905_o ? n1921_o : 1'b0;
  /* decoder.vhd:413:12  */
  assign n1928_o = ~clk_second_cycle_i;
  /* decoder.vhd:414:14  */
  assign n1929_o = ~int_pending_s;
  /* decoder.vhd:414:11  */
  assign n1932_o = n1929_o ? 1'b1 : 1'b0;
  /* decoder.vhd:414:11  */
  assign n1935_o = n1929_o ? 1'b0 : 1'b1;
  /* decoder.vhd:413:9  */
  assign n1937_o = n1928_o ? n1932_o : 1'b0;
  /* decoder.vhd:413:9  */
  assign n1939_o = n1928_o ? n1935_o : 1'b0;
  /* decoder.vhd:397:7  */
  assign n1941_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:422:31  */
  assign n1942_o = ~branch_taken_q;
  /* decoder.vhd:422:27  */
  assign n1943_o = n1942_o & n1905_o;
  /* decoder.vhd:423:12  */
  assign n1944_o = ~int_pending_s;
  /* decoder.vhd:422:50  */
  assign n1945_o = n1944_o & n1943_o;
  /* decoder.vhd:422:9  */
  assign n1948_o = n1945_o ? 1'b1 : 1'b0;
  /* decoder.vhd:421:7  */
  assign n1950_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:428:9  */
  assign n1953_o = n1905_o ? 1'b1 : 1'b0;
  /* decoder.vhd:427:7  */
  assign n1955_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:441:14  */
  assign n1956_o = ~clk_second_cycle_i;
  /* decoder.vhd:441:37  */
  assign n1957_o = assert_psen_s & n1956_o;
  /* decoder.vhd:442:13  */
  assign n1958_o = n1957_o | last_cycle_s;
  /* decoder.vhd:440:23  */
  assign n1959_o = n1958_o & ea_i;
  /* decoder.vhd:440:9  */
  assign n1962_o = n1959_o ? 1'b1 : 1'b0;
  /* decoder.vhd:440:9  */
  assign n1965_o = n1959_o ? 1'b1 : 1'b0;
  /* decoder.vhd:440:9  */
  assign n1968_o = n1959_o ? 1'b1 : 1'b0;
  /* decoder.vhd:439:7  */
  assign n1970_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:450:28  */
  assign n1971_o = n1905_o | last_cycle_s;
  /* decoder.vhd:449:23  */
  assign n1972_o = n1971_o & ea_i;
  /* decoder.vhd:453:12  */
  assign n1973_o = ~p2_output_exp_s;
  /* decoder.vhd:450:45  */
  assign n1974_o = n1973_o & n1972_o;
  /* decoder.vhd:455:12  */
  assign n1975_o = ~movx_first_cycle_s;
  /* decoder.vhd:453:32  */
  assign n1976_o = n1975_o & n1974_o;
  /* decoder.vhd:449:9  */
  assign n1979_o = n1976_o ? 1'b1 : 1'b0;
  /* decoder.vhd:448:7  */
  assign n1981_o = clk_mstate_i == 3'b100;
  assign n1982_o = {n1981_o, n1970_o, n1955_o, n1950_o, n1941_o};
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n1984_o = 1'b0;
      5'b01000: n1984_o = 1'b0;
      5'b00100: n1984_o = 1'b0;
      5'b00010: n1984_o = 1'b0;
      5'b00001: n1984_o = n1923_o;
      default: n1984_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n1987_o = 1'b0;
      5'b01000: n1987_o = n1962_o;
      5'b00100: n1987_o = 1'b0;
      5'b00010: n1987_o = 1'b0;
      5'b00001: n1987_o = 1'b0;
      default: n1987_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n1990_o = 1'b0;
      5'b01000: n1990_o = n1965_o;
      5'b00100: n1990_o = 1'b0;
      5'b00010: n1990_o = 1'b0;
      5'b00001: n1990_o = 1'b0;
      default: n1990_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n1993_o = n1979_o;
      5'b01000: n1993_o = n1968_o;
      5'b00100: n1993_o = 1'b0;
      5'b00010: n1993_o = 1'b0;
      5'b00001: n1993_o = n1925_o;
      default: n1993_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n1996_o = 1'b0;
      5'b01000: n1996_o = 1'b0;
      5'b00100: n1996_o = 1'b0;
      5'b00010: n1996_o = 1'b0;
      5'b00001: n1996_o = n1937_o;
      default: n1996_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n1999_o = 1'b0;
      5'b01000: n1999_o = 1'b0;
      5'b00100: n1999_o = 1'b0;
      5'b00010: n1999_o = 1'b0;
      5'b00001: n1999_o = n1939_o;
      default: n1999_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n2002_o = 1'b0;
      5'b01000: n2002_o = 1'b0;
      5'b00100: n2002_o = 1'b0;
      5'b00010: n2002_o = n1948_o;
      5'b00001: n2002_o = 1'b0;
      default: n2002_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n2005_o = 1'b0;
      5'b01000: n2005_o = 1'b0;
      5'b00100: n2005_o = n1953_o;
      5'b00010: n2005_o = 1'b0;
      5'b00001: n2005_o = 1'b0;
      default: n2005_o = 1'b0;
    endcase
  /* decoder.vhd:396:5  */
  always @*
    case (n1982_o)
      5'b10000: n2008_o = 1'b0;
      5'b01000: n2008_o = 1'b0;
      5'b00100: n2008_o = 1'b0;
      5'b00010: n2008_o = 1'b0;
      5'b00001: n2008_o = n1927_o;
      default: n2008_o = 1'b0;
    endcase
  /* decoder.vhd:615:5  */
  assign n2015_o = int_in_progress_s ? 1'b0 : mb_q;
  /* decoder.vhd:622:8  */
  assign n2016_o = ~clk_second_cycle_i;
  /* decoder.vhd:622:48  */
  assign n2018_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:622:31  */
  assign n2019_o = n2018_o & n2016_o;
  /* decoder.vhd:624:22  */
  assign n2020_o = opc_opcode_q[3];
  /* decoder.vhd:625:43  */
  assign n2021_o = opc_opcode_q[2:0];
  /* decoder.vhd:627:50  */
  assign n2022_o = opc_opcode_q[0];
  /* decoder.vhd:627:36  */
  assign n2024_o = {2'b00, n2022_o};
  /* decoder.vhd:624:7  */
  assign n2025_o = n2020_o ? n2021_o : n2024_o;
  assign n2027_o = n2026_o[7:3];
  /* decoder.vhd:622:5  */
  assign n2030_o = n2019_o ? 1'b1 : 1'b0;
  assign n2032_o = {n2027_o, n2025_o};
  /* decoder.vhd:622:5  */
  assign n2034_o = n2019_o ? n2032_o : 8'bX;
  /* decoder.vhd:622:5  */
  assign n2038_o = n2019_o ? 1'b1 : 1'b0;
  /* decoder.vhd:643:28  */
  assign n2040_o = opc_opcode_q[3];
  /* decoder.vhd:643:32  */
  assign n2041_o = ~n2040_o;
  /* decoder.vhd:642:44  */
  assign n2043_o = 1'b0 | n2041_o;
  /* decoder.vhd:642:13  */
  assign n2050_o = n2043_o ? 1'b1 : n2030_o;
  /* decoder.vhd:642:13  */
  assign n2053_o = n2043_o ? 1'b1 : 1'b0;
  /* decoder.vhd:642:13  */
  assign n2056_o = n2043_o ? 2'b00 : 2'b01;
  /* decoder.vhd:641:11  */
  assign n2058_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:648:11  */
  assign n2063_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:655:28  */
  assign n2067_o = opc_opcode_q[4];
  /* decoder.vhd:655:13  */
  assign n2070_o = n2067_o ? 1'b1 : 1'b0;
  /* decoder.vhd:652:11  */
  assign n2072_o = clk_mstate_i == 3'b100;
  assign n2073_o = {n2072_o, n2063_o, n2058_o};
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2076_o = 1'b1;
      3'b010: n2076_o = 1'b0;
      3'b001: n2076_o = 1'b0;
      default: n2076_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2079_o = 1'b0;
      3'b010: n2079_o = 1'b1;
      3'b001: n2079_o = 1'b0;
      default: n2079_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2082_o = 1'b1;
      3'b010: n2082_o = 1'b0;
      3'b001: n2082_o = 1'b0;
      default: n2082_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2083_o = n2030_o;
      3'b010: n2083_o = n2030_o;
      3'b001: n2083_o = n2050_o;
      default: n2083_o = n2030_o;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2086_o = 1'b0;
      3'b010: n2086_o = 1'b1;
      3'b001: n2086_o = n2053_o;
      default: n2086_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2089_o = 4'b1010;
      3'b010: n2089_o = 4'b1100;
      3'b001: n2089_o = 4'b1100;
      default: n2089_o = 4'b1100;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2091_o = n2070_o;
      3'b010: n2091_o = 1'b0;
      3'b001: n2091_o = 1'b0;
      default: n2091_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2093_o = 2'b01;
      3'b010: n2093_o = 2'b01;
      3'b001: n2093_o = n2056_o;
      default: n2093_o = 2'b01;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2095_o = alu_carry_i;
      3'b010: n2095_o = 1'b0;
      3'b001: n2095_o = 1'b0;
      default: n2095_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2098_o = 1'b1;
      3'b010: n2098_o = 1'b0;
      3'b001: n2098_o = 1'b0;
      default: n2098_o = 1'b0;
    endcase
  /* decoder.vhd:639:9  */
  always @*
    case (n2073_o)
      3'b100: n2101_o = 1'b1;
      3'b010: n2101_o = 1'b0;
      3'b001: n2101_o = 1'b0;
      default: n2101_o = 1'b0;
    endcase
  /* decoder.vhd:638:7  */
  assign n2103_o = opc_mnemonic_s == 6'b000001;
  /* decoder.vhd:675:13  */
  assign n2105_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:682:30  */
  assign n2109_o = opc_opcode_q[4];
  /* decoder.vhd:682:15  */
  assign n2112_o = n2109_o ? 1'b1 : 1'b0;
  /* decoder.vhd:679:13  */
  assign n2114_o = clk_mstate_i == 3'b010;
  assign n2115_o = {n2114_o, n2105_o};
  /* decoder.vhd:673:11  */
  always @*
    case (n2115_o)
      2'b10: n2118_o = 1'b1;
      2'b01: n2118_o = 1'b0;
      default: n2118_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2115_o)
      2'b10: n2121_o = 1'b0;
      2'b01: n2121_o = 1'b1;
      default: n2121_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2115_o)
      2'b10: n2124_o = 1'b1;
      2'b01: n2124_o = 1'b0;
      default: n2124_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2115_o)
      2'b10: n2127_o = 4'b1010;
      2'b01: n2127_o = 4'b1100;
      default: n2127_o = 4'b1100;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2115_o)
      2'b10: n2129_o = n2112_o;
      2'b01: n2129_o = 1'b0;
      default: n2129_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2115_o)
      2'b10: n2131_o = alu_carry_i;
      2'b01: n2131_o = 1'b0;
      default: n2131_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2115_o)
      2'b10: n2134_o = 1'b1;
      2'b01: n2134_o = 1'b0;
      default: n2134_o = 1'b0;
    endcase
  /* decoder.vhd:673:11  */
  always @*
    case (n2115_o)
      2'b10: n2137_o = 1'b1;
      2'b01: n2137_o = 1'b0;
      default: n2137_o = 1'b0;
    endcase
  /* decoder.vhd:672:9  */
  assign n2139_o = clk_second_cycle_i ? n2118_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2141_o = clk_second_cycle_i ? n2121_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2143_o = clk_second_cycle_i ? n2124_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2145_o = clk_second_cycle_i ? n2127_o : 4'b1100;
  /* decoder.vhd:672:9  */
  assign n2147_o = clk_second_cycle_i ? n2129_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2149_o = clk_second_cycle_i ? n2131_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2151_o = clk_second_cycle_i ? n2134_o : 1'b0;
  /* decoder.vhd:672:9  */
  assign n2153_o = clk_second_cycle_i ? n2137_o : 1'b0;
  /* decoder.vhd:669:7  */
  assign n2155_o = opc_mnemonic_s == 6'b000010;
  /* decoder.vhd:703:28  */
  assign n2156_o = opc_opcode_q[3];
  /* decoder.vhd:703:32  */
  assign n2157_o = ~n2156_o;
  /* decoder.vhd:702:44  */
  assign n2159_o = 1'b0 | n2157_o;
  /* decoder.vhd:702:13  */
  assign n2166_o = n2159_o ? 1'b1 : n2030_o;
  /* decoder.vhd:702:13  */
  assign n2169_o = n2159_o ? 1'b1 : 1'b0;
  /* decoder.vhd:702:13  */
  assign n2172_o = n2159_o ? 2'b00 : 2'b01;
  /* decoder.vhd:701:11  */
  assign n2174_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:708:11  */
  assign n2179_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:712:11  */
  assign n2184_o = clk_mstate_i == 3'b100;
  assign n2185_o = {n2184_o, n2179_o, n2174_o};
  /* decoder.vhd:699:9  */
  always @*
    case (n2185_o)
      3'b100: n2188_o = 1'b1;
      3'b010: n2188_o = 1'b0;
      3'b001: n2188_o = 1'b0;
      default: n2188_o = 1'b0;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2185_o)
      3'b100: n2191_o = 1'b0;
      3'b010: n2191_o = 1'b1;
      3'b001: n2191_o = 1'b0;
      default: n2191_o = 1'b0;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2185_o)
      3'b100: n2194_o = 1'b1;
      3'b010: n2194_o = 1'b0;
      3'b001: n2194_o = 1'b0;
      default: n2194_o = 1'b0;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2185_o)
      3'b100: n2195_o = n2030_o;
      3'b010: n2195_o = n2030_o;
      3'b001: n2195_o = n2166_o;
      default: n2195_o = n2030_o;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2185_o)
      3'b100: n2198_o = 1'b0;
      3'b010: n2198_o = 1'b1;
      3'b001: n2198_o = n2169_o;
      default: n2198_o = 1'b0;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2185_o)
      3'b100: n2201_o = 4'b0000;
      3'b010: n2201_o = 4'b1100;
      3'b001: n2201_o = 4'b1100;
      default: n2201_o = 4'b1100;
    endcase
  /* decoder.vhd:699:9  */
  always @*
    case (n2185_o)
      3'b100: n2203_o = 2'b01;
      3'b010: n2203_o = 2'b01;
      3'b001: n2203_o = n2172_o;
      default: n2203_o = 2'b01;
    endcase
  /* decoder.vhd:698:7  */
  assign n2205_o = opc_mnemonic_s == 6'b000011;
  /* decoder.vhd:727:13  */
  assign n2207_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:731:13  */
  assign n2212_o = clk_mstate_i == 3'b010;
  assign n2213_o = {n2212_o, n2207_o};
  /* decoder.vhd:725:11  */
  always @*
    case (n2213_o)
      2'b10: n2216_o = 1'b1;
      2'b01: n2216_o = 1'b0;
      default: n2216_o = 1'b0;
    endcase
  /* decoder.vhd:725:11  */
  always @*
    case (n2213_o)
      2'b10: n2219_o = 1'b0;
      2'b01: n2219_o = 1'b1;
      default: n2219_o = 1'b0;
    endcase
  /* decoder.vhd:725:11  */
  always @*
    case (n2213_o)
      2'b10: n2222_o = 1'b1;
      2'b01: n2222_o = 1'b0;
      default: n2222_o = 1'b0;
    endcase
  /* decoder.vhd:725:11  */
  always @*
    case (n2213_o)
      2'b10: n2225_o = 4'b0000;
      2'b01: n2225_o = 4'b1100;
      default: n2225_o = 4'b1100;
    endcase
  /* decoder.vhd:724:9  */
  assign n2227_o = clk_second_cycle_i ? n2216_o : 1'b0;
  /* decoder.vhd:724:9  */
  assign n2229_o = clk_second_cycle_i ? n2219_o : 1'b0;
  /* decoder.vhd:724:9  */
  assign n2231_o = clk_second_cycle_i ? n2222_o : 1'b0;
  /* decoder.vhd:724:9  */
  assign n2233_o = clk_second_cycle_i ? n2225_o : 4'b1100;
  /* decoder.vhd:721:7  */
  assign n2235_o = opc_mnemonic_s == 6'b000100;
  /* decoder.vhd:745:12  */
  assign n2236_o = ~clk_second_cycle_i;
  /* decoder.vhd:747:27  */
  assign n2238_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:748:28  */
  assign n2239_o = opc_opcode_q[1:0];
  /* decoder.vhd:748:41  */
  assign n2241_o = n2239_o == 2'b00;
  /* decoder.vhd:750:31  */
  assign n2242_o = opc_opcode_q[1];
  /* decoder.vhd:750:35  */
  assign n2243_o = ~n2242_o;
  /* decoder.vhd:750:13  */
  assign n2246_o = n2243_o ? 1'b1 : 1'b0;
  /* decoder.vhd:750:13  */
  assign n2249_o = n2243_o ? 1'b0 : 1'b1;
  /* decoder.vhd:750:13  */
  assign n2252_o = n2243_o ? 1'b1 : 1'b0;
  /* decoder.vhd:750:13  */
  assign n2255_o = n2243_o ? 1'b0 : 1'b1;
  /* decoder.vhd:748:13  */
  assign n2257_o = n2241_o ? 1'b0 : n2246_o;
  /* decoder.vhd:748:13  */
  assign n2259_o = n2241_o ? 1'b0 : n2249_o;
  /* decoder.vhd:748:13  */
  assign n2261_o = n2241_o ? 1'b0 : n2252_o;
  /* decoder.vhd:748:13  */
  assign n2263_o = n2241_o ? 1'b0 : n2255_o;
  /* decoder.vhd:748:13  */
  assign n2266_o = n2241_o ? 1'b1 : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2269_o = n2238_o ? 1'b1 : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2271_o = n2238_o ? n2257_o : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2273_o = n2238_o ? n2259_o : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2275_o = n2238_o ? n2261_o : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2277_o = n2238_o ? n2263_o : 1'b0;
  /* decoder.vhd:747:11  */
  assign n2279_o = n2238_o ? n2266_o : 1'b0;
  /* decoder.vhd:765:13  */
  assign n2281_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:770:13  */
  assign n2283_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:779:30  */
  assign n2284_o = opc_opcode_q[1:0];
  /* decoder.vhd:779:43  */
  assign n2286_o = n2284_o == 2'b00;
  /* decoder.vhd:781:33  */
  assign n2287_o = opc_opcode_q[1];
  /* decoder.vhd:781:37  */
  assign n2288_o = ~n2287_o;
  /* decoder.vhd:781:15  */
  assign n2291_o = n2288_o ? 1'b1 : 1'b0;
  /* decoder.vhd:781:15  */
  assign n2294_o = n2288_o ? 1'b0 : 1'b1;
  /* decoder.vhd:779:15  */
  assign n2297_o = n2286_o ? 1'b1 : 1'b0;
  /* decoder.vhd:779:15  */
  assign n2299_o = n2286_o ? 1'b0 : n2291_o;
  /* decoder.vhd:779:15  */
  assign n2301_o = n2286_o ? 1'b0 : n2294_o;
  /* decoder.vhd:775:13  */
  assign n2303_o = clk_mstate_i == 3'b010;
  assign n2304_o = {n2303_o, n2283_o, n2281_o};
  /* decoder.vhd:762:11  */
  always @*
    case (n2304_o)
      3'b100: n2308_o = 1'b0;
      3'b010: n2308_o = 1'b1;
      3'b001: n2308_o = 1'b1;
      default: n2308_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2304_o)
      3'b100: n2312_o = 1'b1;
      3'b010: n2312_o = 1'b1;
      3'b001: n2312_o = 1'b0;
      default: n2312_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2304_o)
      3'b100: n2314_o = n2297_o;
      3'b010: n2314_o = 1'b0;
      3'b001: n2314_o = 1'b0;
      default: n2314_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2304_o)
      3'b100: n2316_o = n2299_o;
      3'b010: n2316_o = 1'b0;
      3'b001: n2316_o = 1'b0;
      default: n2316_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2304_o)
      3'b100: n2318_o = n2301_o;
      3'b010: n2318_o = 1'b0;
      3'b001: n2318_o = 1'b0;
      default: n2318_o = 1'b0;
    endcase
  /* decoder.vhd:762:11  */
  always @*
    case (n2304_o)
      3'b100: n2321_o = 4'b0000;
      3'b010: n2321_o = 4'b1100;
      3'b001: n2321_o = 4'b1100;
      default: n2321_o = 4'b1100;
    endcase
  /* decoder.vhd:745:9  */
  assign n2323_o = n2236_o ? 1'b0 : n2308_o;
  /* decoder.vhd:745:9  */
  assign n2325_o = n2236_o ? n2269_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2327_o = n2236_o ? 1'b0 : n2312_o;
  /* decoder.vhd:745:9  */
  assign n2329_o = n2236_o ? 1'b0 : n2314_o;
  /* decoder.vhd:745:9  */
  assign n2331_o = n2236_o ? 1'b0 : n2316_o;
  /* decoder.vhd:745:9  */
  assign n2333_o = n2236_o ? n2271_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2335_o = n2236_o ? 1'b0 : n2318_o;
  /* decoder.vhd:745:9  */
  assign n2337_o = n2236_o ? n2273_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2339_o = n2236_o ? 4'b1100 : n2321_o;
  /* decoder.vhd:745:9  */
  assign n2341_o = n2236_o ? n2275_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2343_o = n2236_o ? n2277_o : 1'b0;
  /* decoder.vhd:745:9  */
  assign n2345_o = n2236_o ? n2279_o : 1'b0;
  /* decoder.vhd:742:7  */
  assign n2347_o = opc_mnemonic_s == 6'b000101;
  /* decoder.vhd:798:12  */
  assign n2348_o = ~clk_second_cycle_i;
  /* decoder.vhd:811:18  */
  assign n2349_o = ~int_pending_s;
  /* decoder.vhd:811:15  */
  assign n2352_o = n2349_o ? 1'b1 : 1'b0;
  /* decoder.vhd:802:13  */
  assign n2354_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:816:13  */
  assign n2356_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:822:13  */
  assign n2358_o = clk_mstate_i == 3'b100;
  assign n2359_o = {n2358_o, n2356_o, n2354_o};
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2362_o = 1'b1;
      3'b010: n2362_o = n2030_o;
      3'b001: n2362_o = 1'b1;
      default: n2362_o = n2030_o;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2365_o = 1'b0;
      3'b010: n2365_o = 1'b1;
      3'b001: n2365_o = 1'b0;
      default: n2365_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2368_o = 1'b1;
      3'b010: n2368_o = 1'b0;
      3'b001: n2368_o = 1'b0;
      default: n2368_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2371_o = 1'b1;
      3'b010: n2371_o = 1'b0;
      3'b001: n2371_o = 1'b0;
      default: n2371_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2374_o = 1'b0;
      3'b010: n2374_o = 1'b0;
      3'b001: n2374_o = 1'b1;
      default: n2374_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2378_o = 2'b11;
      3'b010: n2378_o = 2'b01;
      3'b001: n2378_o = 2'b10;
      default: n2378_o = 2'b01;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2381_o = 1'b1;
      3'b010: n2381_o = 1'b0;
      3'b001: n2381_o = 1'b0;
      default: n2381_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2383_o = 1'b0;
      3'b010: n2383_o = 1'b0;
      3'b001: n2383_o = n2352_o;
      default: n2383_o = 1'b0;
    endcase
  /* decoder.vhd:799:11  */
  always @*
    case (n2359_o)
      3'b100: n2387_o = 1'b1;
      3'b010: n2387_o = 1'b1;
      3'b001: n2387_o = 1'b0;
      default: n2387_o = 1'b0;
    endcase
  /* decoder.vhd:845:17  */
  assign n2394_o = tim_int_s ? 1'b0 : 1'b1;
  assign n2395_o = n2389_o[2];
  /* decoder.vhd:845:17  */
  assign n2396_o = tim_int_s ? 1'b1 : n2395_o;
  assign n2397_o = n2389_o[7:3];
  /* decoder.vhd:841:15  */
  assign n2399_o = int_pending_s ? n2394_o : 1'b0;
  assign n2400_o = {n2397_o, n2396_o, 2'b11};
  /* decoder.vhd:841:15  */
  assign n2401_o = int_pending_s ? n2400_o : n2034_o;
  /* decoder.vhd:841:15  */
  assign n2403_o = int_pending_s ? 1'b1 : n2038_o;
  /* decoder.vhd:838:13  */
  assign n2405_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:856:18  */
  assign n2406_o = ~int_pending_s;
  /* decoder.vhd:858:46  */
  assign n2408_o = {4'b0000, n2015_o};
  /* decoder.vhd:858:67  */
  assign n2409_o = opc_opcode_q[7:5];
  /* decoder.vhd:858:53  */
  assign n2410_o = {n2408_o, n2409_o};
  /* decoder.vhd:856:15  */
  assign n2412_o = n2406_o ? n2410_o : 8'b00000000;
  /* decoder.vhd:856:15  */
  assign n2415_o = n2406_o ? 1'b0 : 1'b1;
  /* decoder.vhd:853:13  */
  assign n2417_o = clk_mstate_i == 3'b001;
  assign n2418_o = {n2417_o, n2405_o};
  /* decoder.vhd:836:11  */
  always @*
    case (n2418_o)
      2'b10: n2420_o = 1'b0;
      2'b01: n2420_o = n2399_o;
      default: n2420_o = 1'b0;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2418_o)
      2'b10: n2423_o = 1'b0;
      2'b01: n2423_o = 1'b1;
      default: n2423_o = 1'b0;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2418_o)
      2'b10: n2426_o = 1'b1;
      2'b01: n2426_o = 1'b0;
      default: n2426_o = 1'b0;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2418_o)
      2'b10: n2429_o = 1'b0;
      2'b01: n2429_o = 1'b1;
      default: n2429_o = 1'b0;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2418_o)
      2'b10: n2430_o = n2412_o;
      2'b01: n2430_o = n2401_o;
      default: n2430_o = n2034_o;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2418_o)
      2'b10: n2432_o = 1'b1;
      2'b01: n2432_o = n2403_o;
      default: n2432_o = n2038_o;
    endcase
  /* decoder.vhd:836:11  */
  always @*
    case (n2418_o)
      2'b10: n2434_o = n2415_o;
      2'b01: n2434_o = 1'b0;
      default: n2434_o = 1'b0;
    endcase
  /* decoder.vhd:798:9  */
  assign n2436_o = n2348_o ? 1'b0 : n2420_o;
  /* decoder.vhd:798:9  */
  assign n2437_o = n2348_o ? n2362_o : n2030_o;
  /* decoder.vhd:798:9  */
  assign n2439_o = n2348_o ? 1'b0 : n2423_o;
  /* decoder.vhd:798:9  */
  assign n2441_o = n2348_o ? n2365_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2443_o = n2348_o ? 1'b0 : n2426_o;
  /* decoder.vhd:798:9  */
  assign n2445_o = n2348_o ? n2368_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2447_o = n2348_o ? n2371_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2449_o = n2348_o ? n2374_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2451_o = n2348_o ? n2378_o : 2'b01;
  /* decoder.vhd:798:9  */
  assign n2453_o = n2348_o ? n2381_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2455_o = n2348_o ? 1'b0 : n2429_o;
  /* decoder.vhd:798:9  */
  assign n2457_o = n2348_o ? n2383_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2458_o = n2348_o ? n2034_o : n2430_o;
  /* decoder.vhd:798:9  */
  assign n2459_o = n2348_o ? n2038_o : n2432_o;
  /* decoder.vhd:798:9  */
  assign n2461_o = n2348_o ? n2387_o : 1'b0;
  /* decoder.vhd:798:9  */
  assign n2463_o = n2348_o ? 1'b0 : n2434_o;
  /* decoder.vhd:795:7  */
  assign n2465_o = opc_mnemonic_s == 6'b000110;
  /* decoder.vhd:875:25  */
  assign n2467_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:875:9  */
  assign n2470_o = n2467_o ? 1'b1 : 1'b0;
  /* decoder.vhd:875:9  */
  assign n2473_o = n2467_o ? 1'b1 : 1'b0;
  /* decoder.vhd:875:9  */
  assign n2476_o = n2467_o ? 4'b0100 : 4'b1100;
  /* decoder.vhd:873:7  */
  assign n2478_o = opc_mnemonic_s == 6'b000111;
  /* decoder.vhd:884:25  */
  assign n2480_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:884:9  */
  assign n2483_o = n2480_o ? 1'b1 : 1'b0;
  /* decoder.vhd:882:7  */
  assign n2485_o = opc_mnemonic_s == 6'b001000;
  /* decoder.vhd:892:25  */
  assign n2487_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:893:26  */
  assign n2488_o = opc_opcode_q[5];
  /* decoder.vhd:893:30  */
  assign n2489_o = ~n2488_o;
  /* decoder.vhd:893:11  */
  assign n2492_o = n2489_o ? 1'b1 : 1'b0;
  /* decoder.vhd:893:11  */
  assign n2495_o = n2489_o ? 1'b0 : 1'b1;
  /* decoder.vhd:892:9  */
  assign n2497_o = n2487_o ? n2492_o : 1'b0;
  /* decoder.vhd:892:9  */
  assign n2499_o = n2487_o ? n2495_o : 1'b0;
  /* decoder.vhd:890:7  */
  assign n2501_o = opc_mnemonic_s == 6'b001001;
  /* decoder.vhd:905:25  */
  assign n2503_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:905:9  */
  assign n2506_o = n2503_o ? 1'b1 : 1'b0;
  /* decoder.vhd:905:9  */
  assign n2509_o = n2503_o ? 1'b1 : 1'b0;
  /* decoder.vhd:905:9  */
  assign n2512_o = n2503_o ? 4'b0011 : 4'b1100;
  /* decoder.vhd:903:7  */
  assign n2514_o = opc_mnemonic_s == 6'b001010;
  /* decoder.vhd:914:25  */
  assign n2516_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:915:33  */
  assign n2517_o = ~psw_carry_i;
  /* decoder.vhd:914:9  */
  assign n2519_o = n2516_o ? n2517_o : 1'b0;
  /* decoder.vhd:914:9  */
  assign n2522_o = n2516_o ? 1'b1 : 1'b0;
  /* decoder.vhd:912:7  */
  assign n2524_o = opc_mnemonic_s == 6'b001011;
  /* decoder.vhd:922:25  */
  assign n2526_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:923:26  */
  assign n2527_o = opc_opcode_q[5];
  /* decoder.vhd:923:30  */
  assign n2528_o = ~n2527_o;
  /* decoder.vhd:924:35  */
  assign n2529_o = ~psw_f0_i;
  /* decoder.vhd:923:11  */
  assign n2531_o = n2528_o ? n2529_o : 1'b0;
  /* decoder.vhd:923:11  */
  assign n2534_o = n2528_o ? 1'b1 : 1'b0;
  /* decoder.vhd:923:11  */
  assign n2537_o = n2528_o ? 1'b0 : 1'b1;
  /* decoder.vhd:922:9  */
  assign n2539_o = n2526_o ? n2531_o : 1'b0;
  /* decoder.vhd:922:9  */
  assign n2541_o = n2526_o ? n2534_o : 1'b0;
  /* decoder.vhd:922:9  */
  assign n2543_o = n2526_o ? n2537_o : 1'b0;
  /* decoder.vhd:920:7  */
  assign n2545_o = opc_mnemonic_s == 6'b001100;
  /* decoder.vhd:938:11  */
  assign n2547_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:944:38  */
  assign n2548_o = psw_aux_carry_i | alu_da_overflow_i;
  /* decoder.vhd:944:13  */
  assign n2551_o = n2548_o ? 1'b1 : 1'b0;
  /* decoder.vhd:944:13  */
  assign n2554_o = n2548_o ? 1'b1 : 1'b0;
  /* decoder.vhd:943:11  */
  assign n2556_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:958:13  */
  assign n2559_o = alu_da_overflow_i ? 4'b1010 : 4'b1100;
  /* decoder.vhd:958:13  */
  assign n2561_o = alu_da_overflow_i ? alu_carry_i : 1'b0;
  /* decoder.vhd:955:11  */
  assign n2563_o = clk_mstate_i == 3'b100;
  assign n2564_o = {n2563_o, n2556_o, n2547_o};
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2567_o = 1'b1;
      3'b010: n2567_o = 1'b0;
      3'b001: n2567_o = 1'b0;
      default: n2567_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2569_o = 1'b0;
      3'b010: n2569_o = n2551_o;
      3'b001: n2569_o = 1'b0;
      default: n2569_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2572_o = 1'b1;
      3'b010: n2572_o = n2554_o;
      3'b001: n2572_o = 1'b0;
      default: n2572_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2574_o = n2559_o;
      3'b010: n2574_o = 4'b1010;
      3'b001: n2574_o = 4'b1010;
      default: n2574_o = 4'b1010;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2578_o = 1'b1;
      3'b010: n2578_o = 1'b0;
      3'b001: n2578_o = 1'b0;
      default: n2578_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2581_o = 1'b0;
      3'b010: n2581_o = 1'b0;
      3'b001: n2581_o = 1'b1;
      default: n2581_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2584_o = 1'b0;
      3'b010: n2584_o = 1'b1;
      3'b001: n2584_o = 1'b0;
      default: n2584_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2586_o = n2561_o;
      3'b010: n2586_o = 1'b0;
      3'b001: n2586_o = 1'b0;
      default: n2586_o = 1'b0;
    endcase
  /* decoder.vhd:936:9  */
  always @*
    case (n2564_o)
      3'b100: n2589_o = 1'b1;
      3'b010: n2589_o = 1'b0;
      3'b001: n2589_o = 1'b0;
      default: n2589_o = 1'b0;
    endcase
  /* decoder.vhd:933:7  */
  assign n2591_o = opc_mnemonic_s == 6'b001101;
  /* decoder.vhd:978:28  */
  assign n2592_o = opc_opcode_q[6];
  /* decoder.vhd:978:13  */
  assign n2595_o = n2592_o ? 1'b1 : 1'b0;
  /* decoder.vhd:978:13  */
  assign n2598_o = n2592_o ? 1'b1 : 1'b0;
  /* decoder.vhd:976:11  */
  assign n2600_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:987:28  */
  assign n2601_o = opc_opcode_q[6];
  /* decoder.vhd:987:32  */
  assign n2602_o = ~n2601_o;
  /* decoder.vhd:987:13  */
  assign n2605_o = n2602_o ? 1'b1 : 1'b0;
  /* decoder.vhd:987:13  */
  assign n2608_o = n2602_o ? 1'b0 : 1'b1;
  /* decoder.vhd:983:11  */
  assign n2610_o = clk_mstate_i == 3'b100;
  assign n2611_o = {n2610_o, n2600_o};
  /* decoder.vhd:975:9  */
  always @*
    case (n2611_o)
      2'b10: n2613_o = n2605_o;
      2'b01: n2613_o = 1'b0;
      default: n2613_o = 1'b0;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2611_o)
      2'b10: n2615_o = 1'b0;
      2'b01: n2615_o = n2595_o;
      default: n2615_o = 1'b0;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2611_o)
      2'b10: n2618_o = 1'b1;
      2'b01: n2618_o = 1'b0;
      default: n2618_o = 1'b0;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2611_o)
      2'b10: n2620_o = 1'b0;
      2'b01: n2620_o = n2598_o;
      default: n2620_o = 1'b0;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2611_o)
      2'b10: n2623_o = 4'b1000;
      2'b01: n2623_o = 4'b1100;
      default: n2623_o = 4'b1100;
    endcase
  /* decoder.vhd:975:9  */
  always @*
    case (n2611_o)
      2'b10: n2625_o = n2608_o;
      2'b01: n2625_o = 1'b0;
      default: n2625_o = 1'b0;
    endcase
  /* decoder.vhd:974:7  */
  assign n2627_o = opc_mnemonic_s == 6'b001110;
  /* decoder.vhd:1002:25  */
  assign n2629_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1003:26  */
  assign n2630_o = opc_opcode_q[4];
  /* decoder.vhd:1003:11  */
  assign n2633_o = n2630_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1003:11  */
  assign n2636_o = n2630_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1002:9  */
  assign n2638_o = n2629_o ? n2633_o : 1'b0;
  /* decoder.vhd:1002:9  */
  assign n2640_o = n2629_o ? n2636_o : 1'b0;
  /* decoder.vhd:1001:7  */
  assign n2642_o = opc_mnemonic_s == 6'b001111;
  /* decoder.vhd:1012:25  */
  assign n2644_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1013:26  */
  assign n2645_o = opc_opcode_q[4];
  /* decoder.vhd:1013:11  */
  assign n2648_o = n2645_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1013:11  */
  assign n2651_o = n2645_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1012:9  */
  assign n2653_o = n2644_o ? n2648_o : 1'b0;
  /* decoder.vhd:1012:9  */
  assign n2655_o = n2644_o ? n2651_o : 1'b0;
  /* decoder.vhd:1011:7  */
  assign n2657_o = opc_mnemonic_s == 6'b010000;
  /* decoder.vhd:1024:12  */
  assign n2658_o = ~clk_second_cycle_i;
  /* decoder.vhd:1027:13  */
  assign n2660_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1033:13  */
  assign n2663_o = clk_mstate_i == 3'b100;
  assign n2664_o = {n2663_o, n2660_o};
  /* decoder.vhd:1025:11  */
  always @*
    case (n2664_o)
      2'b10: n2667_o = 1'b0;
      2'b01: n2667_o = 1'b1;
      default: n2667_o = 1'b0;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2664_o)
      2'b10: n2670_o = 1'b1;
      2'b01: n2670_o = 1'b0;
      default: n2670_o = 1'b0;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2664_o)
      2'b10: n2673_o = 1'b0;
      2'b01: n2673_o = 1'b1;
      default: n2673_o = 1'b0;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2664_o)
      2'b10: n2676_o = 4'b1000;
      2'b01: n2676_o = 4'b1100;
      default: n2676_o = 4'b1100;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2664_o)
      2'b10: n2679_o = 1'b1;
      2'b01: n2679_o = 1'b0;
      default: n2679_o = 1'b0;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2664_o)
      2'b10: n2682_o = 4'b0001;
      2'b01: n2682_o = 4'b0000;
      default: n2682_o = 4'b0000;
    endcase
  assign n2683_o = opc_opcode_q[5];
  /* decoder.vhd:1025:11  */
  always @*
    case (n2664_o)
      2'b10: n2684_o = 1'b0;
      2'b01: n2684_o = n2683_o;
      default: n2684_o = n2683_o;
    endcase
  /* decoder.vhd:1025:11  */
  always @*
    case (n2664_o)
      2'b10: n2687_o = 1'b1;
      2'b01: n2687_o = 1'b0;
      default: n2687_o = 1'b0;
    endcase
  /* decoder.vhd:1050:27  */
  assign n2689_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1050:37  */
  assign n2690_o = cnd_take_branch_i & n2689_o;
  /* decoder.vhd:1050:11  */
  assign n2696_o = n2690_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1050:11  */
  assign n2699_o = n2690_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2701_o = n2658_o ? n2667_o : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2703_o = n2658_o ? n2670_o : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2705_o = n2658_o ? n2673_o : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2707_o = n2658_o ? 1'b0 : n2696_o;
  /* decoder.vhd:1024:9  */
  assign n2709_o = n2658_o ? n2676_o : 4'b1100;
  /* decoder.vhd:1024:9  */
  assign n2711_o = n2658_o ? n2679_o : 1'b0;
  /* decoder.vhd:1024:9  */
  assign n2713_o = n2658_o ? n2682_o : 4'b0000;
  assign n2714_o = opc_opcode_q[5];
  /* decoder.vhd:1024:9  */
  assign n2715_o = n2658_o ? n2684_o : n2714_o;
  /* decoder.vhd:1024:9  */
  assign n2717_o = n2658_o ? 1'b0 : n2699_o;
  /* decoder.vhd:1024:9  */
  assign n2719_o = n2658_o ? n2687_o : 1'b0;
  /* decoder.vhd:1021:7  */
  assign n2721_o = opc_mnemonic_s == 6'b010001;
  /* decoder.vhd:1058:25  */
  assign n2723_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1059:26  */
  assign n2724_o = opc_opcode_q[4];
  /* decoder.vhd:1059:30  */
  assign n2725_o = ~n2724_o;
  /* decoder.vhd:1059:11  */
  assign n2728_o = n2725_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1059:11  */
  assign n2731_o = n2725_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1058:9  */
  assign n2733_o = n2723_o ? n2728_o : 1'b0;
  /* decoder.vhd:1058:9  */
  assign n2735_o = n2723_o ? n2731_o : 1'b0;
  /* decoder.vhd:1057:7  */
  assign n2737_o = opc_mnemonic_s == 6'b111110;
  /* decoder.vhd:1068:25  */
  assign n2739_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1068:9  */
  assign n2742_o = n2739_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1067:7  */
  assign n2744_o = opc_mnemonic_s == 6'b010010;
  /* decoder.vhd:1075:48  */
  assign n2746_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1075:31  */
  assign n2747_o = n2746_o & clk_second_cycle_i;
  /* decoder.vhd:1078:26  */
  assign n2748_o = opc_opcode_q[1];
  /* decoder.vhd:1078:30  */
  assign n2749_o = ~n2748_o;
  /* decoder.vhd:1078:11  */
  assign n2752_o = n2749_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1078:11  */
  assign n2755_o = n2749_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1075:9  */
  assign n2758_o = n2747_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1075:9  */
  assign n2760_o = n2747_o ? n2752_o : 1'b0;
  /* decoder.vhd:1075:9  */
  assign n2762_o = n2747_o ? n2755_o : 1'b0;
  /* decoder.vhd:1073:7  */
  assign n2764_o = opc_mnemonic_s == 6'b010011;
  /* decoder.vhd:1088:25  */
  assign n2766_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1088:9  */
  assign n2769_o = n2766_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1088:9  */
  assign n2772_o = n2766_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1086:7  */
  assign n2774_o = opc_mnemonic_s == 6'b111010;
  /* decoder.vhd:1099:48  */
  assign n2776_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1099:31  */
  assign n2777_o = n2776_o & clk_second_cycle_i;
  /* decoder.vhd:1099:9  */
  assign n2780_o = n2777_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1099:9  */
  assign n2783_o = n2777_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1095:7  */
  assign n2785_o = opc_mnemonic_s == 6'b010101;
  /* decoder.vhd:1111:28  */
  assign n2786_o = opc_opcode_q[3];
  /* decoder.vhd:1111:32  */
  assign n2787_o = ~n2786_o;
  /* decoder.vhd:1110:44  */
  assign n2789_o = 1'b0 | n2787_o;
  /* decoder.vhd:1110:13  */
  assign n2796_o = n2789_o ? 1'b1 : n2030_o;
  /* decoder.vhd:1110:13  */
  assign n2799_o = n2789_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1110:13  */
  assign n2802_o = n2789_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1109:11  */
  assign n2804_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1117:28  */
  assign n2805_o = opc_opcode_q[3:2];
  /* decoder.vhd:1117:41  */
  assign n2807_o = n2805_o != 2'b01;
  /* decoder.vhd:1117:13  */
  assign n2810_o = n2807_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1117:13  */
  assign n2813_o = n2807_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1115:11  */
  assign n2815_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1126:28  */
  assign n2816_o = opc_opcode_q[3:2];
  /* decoder.vhd:1126:41  */
  assign n2818_o = n2816_o == 2'b01;
  /* decoder.vhd:1126:13  */
  assign n2821_o = n2818_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1126:13  */
  assign n2824_o = n2818_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1122:11  */
  assign n2826_o = clk_mstate_i == 3'b100;
  assign n2827_o = {n2826_o, n2815_o, n2804_o};
  /* decoder.vhd:1107:9  */
  always @*
    case (n2827_o)
      3'b100: n2829_o = n2821_o;
      3'b010: n2829_o = 1'b0;
      3'b001: n2829_o = 1'b0;
      default: n2829_o = 1'b0;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2827_o)
      3'b100: n2831_o = 1'b0;
      3'b010: n2831_o = n2810_o;
      3'b001: n2831_o = 1'b0;
      default: n2831_o = 1'b0;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2827_o)
      3'b100: n2834_o = 1'b1;
      3'b010: n2834_o = 1'b0;
      3'b001: n2834_o = 1'b0;
      default: n2834_o = 1'b0;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2827_o)
      3'b100: n2835_o = n2030_o;
      3'b010: n2835_o = n2030_o;
      3'b001: n2835_o = n2796_o;
      default: n2835_o = n2030_o;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2827_o)
      3'b100: n2837_o = 1'b0;
      3'b010: n2837_o = n2813_o;
      3'b001: n2837_o = n2799_o;
      default: n2837_o = 1'b0;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2827_o)
      3'b100: n2840_o = 4'b1001;
      3'b010: n2840_o = 4'b1100;
      3'b001: n2840_o = 4'b1100;
      default: n2840_o = 4'b1100;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2827_o)
      3'b100: n2842_o = 2'b01;
      3'b010: n2842_o = 2'b01;
      3'b001: n2842_o = n2802_o;
      default: n2842_o = 2'b01;
    endcase
  /* decoder.vhd:1107:9  */
  always @*
    case (n2827_o)
      3'b100: n2844_o = n2824_o;
      3'b010: n2844_o = 1'b0;
      3'b001: n2844_o = 1'b0;
      default: n2844_o = 1'b0;
    endcase
  /* decoder.vhd:1106:7  */
  assign n2846_o = opc_mnemonic_s == 6'b010100;
  /* decoder.vhd:1144:12  */
  assign n2847_o = ~clk_second_cycle_i;
  /* decoder.vhd:1146:27  */
  assign n2849_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1146:11  */
  assign n2852_o = n2849_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1146:11  */
  assign n2855_o = n2849_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1155:27  */
  assign n2857_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1155:37  */
  assign n2858_o = cnd_take_branch_i & n2857_o;
  /* decoder.vhd:1155:11  */
  assign n2864_o = n2858_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1155:11  */
  assign n2867_o = n2858_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1144:9  */
  assign n2869_o = n2847_o ? n2852_o : 1'b0;
  /* decoder.vhd:1144:9  */
  assign n2871_o = n2847_o ? 1'b0 : n2864_o;
  /* decoder.vhd:1144:9  */
  assign n2873_o = n2847_o ? n2855_o : 1'b0;
  /* decoder.vhd:1144:9  */
  assign n2875_o = n2847_o ? 1'b0 : n2867_o;
  /* decoder.vhd:1140:7  */
  assign n2877_o = opc_mnemonic_s == 6'b010110;
  /* decoder.vhd:1166:12  */
  assign n2878_o = ~clk_second_cycle_i;
  /* decoder.vhd:1168:27  */
  assign n2880_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1170:48  */
  assign n2881_o = opc_opcode_q[4];
  /* decoder.vhd:1168:11  */
  assign n2884_o = n2880_o ? 1'b1 : 1'b0;
  assign n2885_o = opc_opcode_q[5];
  /* decoder.vhd:1166:9  */
  assign n2886_o = n2904_o ? n2881_o : n2885_o;
  /* decoder.vhd:1176:27  */
  assign n2888_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1176:37  */
  assign n2889_o = cnd_take_branch_i & n2888_o;
  /* decoder.vhd:1176:11  */
  assign n2895_o = n2889_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1176:11  */
  assign n2898_o = n2889_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1166:9  */
  assign n2900_o = n2878_o ? 1'b0 : n2895_o;
  /* decoder.vhd:1166:9  */
  assign n2902_o = n2878_o ? n2884_o : 1'b0;
  /* decoder.vhd:1166:9  */
  assign n2904_o = n2878_o & n2880_o;
  /* decoder.vhd:1166:9  */
  assign n2906_o = n2878_o ? 1'b0 : n2898_o;
  /* decoder.vhd:1162:7  */
  assign n2908_o = opc_mnemonic_s == 6'b010111;
  /* decoder.vhd:1186:12  */
  assign n2909_o = ~clk_second_cycle_i;
  /* decoder.vhd:1188:27  */
  assign n2911_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1190:28  */
  assign n2912_o = opc_opcode_q[7];
  /* decoder.vhd:1190:13  */
  assign n2915_o = n2912_o ? 4'b0011 : 4'b0100;
  /* decoder.vhd:1188:11  */
  assign n2918_o = n2911_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1188:11  */
  assign n2920_o = n2911_o ? n2915_o : 4'b0000;
  /* decoder.vhd:1203:27  */
  assign n2922_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1203:37  */
  assign n2923_o = cnd_take_branch_i & n2922_o;
  /* decoder.vhd:1203:11  */
  assign n2929_o = n2923_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1203:11  */
  assign n2932_o = n2923_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1186:9  */
  assign n2934_o = n2909_o ? 1'b0 : n2929_o;
  /* decoder.vhd:1186:9  */
  assign n2936_o = n2909_o ? n2918_o : 1'b0;
  /* decoder.vhd:1186:9  */
  assign n2938_o = n2909_o ? n2920_o : 4'b0000;
  /* decoder.vhd:1186:9  */
  assign n2940_o = n2909_o ? 1'b0 : n2932_o;
  /* decoder.vhd:1183:7  */
  assign n2942_o = opc_mnemonic_s == 6'b011000;
  /* decoder.vhd:1217:13  */
  assign n2944_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1223:40  */
  assign n2946_o = {4'b0000, n2015_o};
  /* decoder.vhd:1223:61  */
  assign n2947_o = opc_opcode_q[7:5];
  /* decoder.vhd:1223:47  */
  assign n2948_o = {n2946_o, n2947_o};
  /* decoder.vhd:1222:13  */
  assign n2950_o = clk_mstate_i == 3'b001;
  assign n2951_o = {n2950_o, n2944_o};
  /* decoder.vhd:1215:11  */
  always @*
    case (n2951_o)
      2'b10: n2954_o = 1'b0;
      2'b01: n2954_o = 1'b1;
      default: n2954_o = 1'b0;
    endcase
  /* decoder.vhd:1215:11  */
  always @*
    case (n2951_o)
      2'b10: n2957_o = 1'b1;
      2'b01: n2957_o = 1'b0;
      default: n2957_o = 1'b0;
    endcase
  /* decoder.vhd:1215:11  */
  always @*
    case (n2951_o)
      2'b10: n2960_o = 1'b0;
      2'b01: n2960_o = 1'b1;
      default: n2960_o = 1'b0;
    endcase
  /* decoder.vhd:1215:11  */
  always @*
    case (n2951_o)
      2'b10: n2961_o = n2948_o;
      2'b01: n2961_o = n2034_o;
      default: n2961_o = n2034_o;
    endcase
  /* decoder.vhd:1215:11  */
  always @*
    case (n2951_o)
      2'b10: n2963_o = 1'b1;
      2'b01: n2963_o = n2038_o;
      default: n2963_o = n2038_o;
    endcase
  /* decoder.vhd:1214:9  */
  assign n2965_o = clk_second_cycle_i ? n2954_o : 1'b0;
  /* decoder.vhd:1214:9  */
  assign n2967_o = clk_second_cycle_i ? n2957_o : 1'b0;
  /* decoder.vhd:1214:9  */
  assign n2969_o = clk_second_cycle_i ? n2960_o : 1'b0;
  /* decoder.vhd:1214:9  */
  assign n2970_o = clk_second_cycle_i ? n2961_o : n2034_o;
  /* decoder.vhd:1214:9  */
  assign n2971_o = clk_second_cycle_i ? n2963_o : n2038_o;
  /* decoder.vhd:1211:7  */
  assign n2973_o = opc_mnemonic_s == 6'b011001;
  /* decoder.vhd:1238:12  */
  assign n2974_o = ~clk_second_cycle_i;
  /* decoder.vhd:1241:27  */
  assign n2976_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1241:11  */
  assign n2979_o = n2976_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1241:11  */
  assign n2982_o = n2976_o ? 2'b01 : 2'b00;
  /* decoder.vhd:1247:27  */
  assign n2984_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1247:11  */
  assign n2987_o = n2984_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1247:11  */
  assign n2990_o = n2984_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1238:9  */
  assign n2992_o = n2974_o ? n2979_o : 1'b0;
  /* decoder.vhd:1238:9  */
  assign n2994_o = n2974_o ? 1'b0 : n2987_o;
  /* decoder.vhd:1238:9  */
  assign n2996_o = n2974_o ? n2982_o : 2'b00;
  /* decoder.vhd:1238:9  */
  assign n2998_o = n2974_o ? 1'b0 : n2990_o;
  /* decoder.vhd:1235:7  */
  assign n3000_o = opc_mnemonic_s == 6'b011010;
  /* decoder.vhd:1260:12  */
  assign n3001_o = ~clk_second_cycle_i;
  /* decoder.vhd:1262:27  */
  assign n3003_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1262:11  */
  assign n3006_o = n3003_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1269:27  */
  assign n3008_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1269:37  */
  assign n3009_o = cnd_take_branch_i & n3008_o;
  /* decoder.vhd:1269:11  */
  assign n3015_o = n3009_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1269:11  */
  assign n3018_o = n3009_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1260:9  */
  assign n3020_o = n3001_o ? 1'b0 : n3015_o;
  /* decoder.vhd:1260:9  */
  assign n3022_o = n3001_o ? n3006_o : 1'b0;
  /* decoder.vhd:1260:9  */
  assign n3024_o = n3001_o ? 1'b0 : n3018_o;
  /* decoder.vhd:1256:7  */
  assign n3026_o = opc_mnemonic_s == 6'b011011;
  /* decoder.vhd:1280:12  */
  assign n3027_o = ~clk_second_cycle_i;
  /* decoder.vhd:1282:27  */
  assign n3029_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1282:11  */
  assign n3032_o = n3029_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1289:27  */
  assign n3034_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1289:37  */
  assign n3035_o = cnd_take_branch_i & n3034_o;
  /* decoder.vhd:1289:11  */
  assign n3041_o = n3035_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1289:11  */
  assign n3044_o = n3035_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1280:9  */
  assign n3046_o = n3027_o ? 1'b0 : n3041_o;
  /* decoder.vhd:1280:9  */
  assign n3048_o = n3027_o ? n3032_o : 1'b0;
  /* decoder.vhd:1280:9  */
  assign n3050_o = n3027_o ? 1'b0 : n3044_o;
  /* decoder.vhd:1276:7  */
  assign n3052_o = opc_mnemonic_s == 6'b111100;
  /* decoder.vhd:1300:12  */
  assign n3053_o = ~clk_second_cycle_i;
  /* decoder.vhd:1302:27  */
  assign n3055_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1302:11  */
  assign n3058_o = n3055_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1309:27  */
  assign n3060_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1309:37  */
  assign n3061_o = cnd_take_branch_i & n3060_o;
  /* decoder.vhd:1309:11  */
  assign n3067_o = n3061_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1309:11  */
  assign n3070_o = n3061_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1300:9  */
  assign n3072_o = n3053_o ? 1'b0 : n3067_o;
  /* decoder.vhd:1300:9  */
  assign n3074_o = n3053_o ? n3058_o : 1'b0;
  /* decoder.vhd:1300:9  */
  assign n3076_o = n3053_o ? 1'b0 : n3070_o;
  /* decoder.vhd:1296:7  */
  assign n3078_o = opc_mnemonic_s == 6'b111101;
  /* decoder.vhd:1318:24  */
  assign n3079_o = opc_opcode_q[6];
  /* decoder.vhd:1318:28  */
  assign n3080_o = ~n3079_o;
  /* decoder.vhd:1318:9  */
  assign n3083_o = n3080_o ? 4'b0110 : 4'b0111;
  /* decoder.vhd:1324:12  */
  assign n3084_o = ~clk_second_cycle_i;
  /* decoder.vhd:1326:27  */
  assign n3086_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1328:48  */
  assign n3087_o = opc_opcode_q[4];
  /* decoder.vhd:1326:11  */
  assign n3090_o = n3086_o ? 1'b1 : 1'b0;
  assign n3091_o = opc_opcode_q[5];
  /* decoder.vhd:1324:9  */
  assign n3092_o = n3110_o ? n3087_o : n3091_o;
  /* decoder.vhd:1334:27  */
  assign n3094_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1334:37  */
  assign n3095_o = cnd_take_branch_i & n3094_o;
  /* decoder.vhd:1334:11  */
  assign n3101_o = n3095_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1334:11  */
  assign n3104_o = n3095_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1324:9  */
  assign n3106_o = n3084_o ? 1'b0 : n3101_o;
  /* decoder.vhd:1324:9  */
  assign n3108_o = n3084_o ? n3090_o : 1'b0;
  /* decoder.vhd:1324:9  */
  assign n3110_o = n3084_o & n3086_o;
  /* decoder.vhd:1324:9  */
  assign n3112_o = n3084_o ? 1'b0 : n3104_o;
  /* decoder.vhd:1316:7  */
  assign n3114_o = opc_mnemonic_s == 6'b011100;
  /* decoder.vhd:1345:12  */
  assign n3115_o = ~clk_second_cycle_i;
  /* decoder.vhd:1347:27  */
  assign n3117_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1347:11  */
  assign n3120_o = n3117_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1347:11  */
  assign n3123_o = n3117_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1355:27  */
  assign n3125_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1355:37  */
  assign n3126_o = cnd_take_branch_i & n3125_o;
  /* decoder.vhd:1355:11  */
  assign n3132_o = n3126_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1355:11  */
  assign n3135_o = n3126_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1345:9  */
  assign n3137_o = n3115_o ? 1'b0 : n3132_o;
  /* decoder.vhd:1345:9  */
  assign n3139_o = n3115_o ? n3120_o : 1'b0;
  /* decoder.vhd:1345:9  */
  assign n3141_o = n3115_o ? 1'b0 : n3135_o;
  /* decoder.vhd:1345:9  */
  assign n3143_o = n3115_o ? n3123_o : 1'b0;
  /* decoder.vhd:1341:7  */
  assign n3145_o = opc_mnemonic_s == 6'b011101;
  /* decoder.vhd:1366:12  */
  assign n3146_o = ~clk_second_cycle_i;
  /* decoder.vhd:1368:27  */
  assign n3148_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1371:48  */
  assign n3149_o = opc_opcode_q[6];
  /* decoder.vhd:1368:11  */
  assign n3152_o = n3148_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1368:11  */
  assign n3155_o = n3148_o ? 1'b1 : 1'b0;
  assign n3156_o = opc_opcode_q[5];
  /* decoder.vhd:1366:9  */
  assign n3157_o = n3177_o ? n3149_o : n3156_o;
  /* decoder.vhd:1377:27  */
  assign n3159_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1377:37  */
  assign n3160_o = cnd_take_branch_i & n3159_o;
  /* decoder.vhd:1377:11  */
  assign n3166_o = n3160_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1377:11  */
  assign n3169_o = n3160_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1366:9  */
  assign n3171_o = n3146_o ? n3152_o : 1'b0;
  /* decoder.vhd:1366:9  */
  assign n3173_o = n3146_o ? 1'b0 : n3166_o;
  /* decoder.vhd:1366:9  */
  assign n3175_o = n3146_o ? n3155_o : 1'b0;
  /* decoder.vhd:1366:9  */
  assign n3177_o = n3146_o & n3148_o;
  /* decoder.vhd:1366:9  */
  assign n3179_o = n3146_o ? 1'b0 : n3169_o;
  /* decoder.vhd:1362:7  */
  assign n3181_o = opc_mnemonic_s == 6'b011110;
  /* decoder.vhd:1389:48  */
  assign n3183_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1389:31  */
  assign n3184_o = n3183_o & clk_second_cycle_i;
  /* decoder.vhd:1389:9  */
  assign n3187_o = n3184_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1384:7  */
  assign n3189_o = opc_mnemonic_s == 6'b011111;
  /* decoder.vhd:1399:28  */
  assign n3190_o = opc_opcode_q[3];
  /* decoder.vhd:1399:32  */
  assign n3191_o = ~n3190_o;
  /* decoder.vhd:1398:44  */
  assign n3193_o = 1'b0 | n3191_o;
  /* decoder.vhd:1398:13  */
  assign n3200_o = n3193_o ? 1'b1 : n2030_o;
  /* decoder.vhd:1398:13  */
  assign n3203_o = n3193_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1398:13  */
  assign n3206_o = n3193_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1397:11  */
  assign n3208_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1404:11  */
  assign n3213_o = clk_mstate_i == 3'b011;
  assign n3214_o = {n3213_o, n3208_o};
  /* decoder.vhd:1395:9  */
  always @*
    case (n3214_o)
      2'b10: n3217_o = 1'b1;
      2'b01: n3217_o = 1'b0;
      default: n3217_o = 1'b0;
    endcase
  /* decoder.vhd:1395:9  */
  always @*
    case (n3214_o)
      2'b10: n3220_o = 1'b1;
      2'b01: n3220_o = 1'b0;
      default: n3220_o = 1'b0;
    endcase
  /* decoder.vhd:1395:9  */
  always @*
    case (n3214_o)
      2'b10: n3221_o = n2030_o;
      2'b01: n3221_o = n3200_o;
      default: n3221_o = n2030_o;
    endcase
  /* decoder.vhd:1395:9  */
  always @*
    case (n3214_o)
      2'b10: n3224_o = 1'b1;
      2'b01: n3224_o = n3203_o;
      default: n3224_o = 1'b0;
    endcase
  /* decoder.vhd:1395:9  */
  always @*
    case (n3214_o)
      2'b10: n3226_o = 2'b01;
      2'b01: n3226_o = n3206_o;
      default: n3226_o = 2'b01;
    endcase
  /* decoder.vhd:1394:7  */
  assign n3228_o = opc_mnemonic_s == 6'b100001;
  /* decoder.vhd:1415:25  */
  assign n3230_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1415:9  */
  assign n3233_o = n3230_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1415:9  */
  assign n3236_o = n3230_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1415:9  */
  assign n3239_o = n3230_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1414:7  */
  assign n3241_o = opc_mnemonic_s == 6'b100000;
  /* decoder.vhd:1423:25  */
  assign n3243_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1423:9  */
  assign n3246_o = n3243_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1423:9  */
  assign n3249_o = n3243_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1423:9  */
  assign n3252_o = n3243_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1422:7  */
  assign n3254_o = opc_mnemonic_s == 6'b100010;
  /* decoder.vhd:1435:28  */
  assign n3255_o = opc_opcode_q[3];
  /* decoder.vhd:1435:32  */
  assign n3256_o = ~n3255_o;
  /* decoder.vhd:1434:44  */
  assign n3258_o = 1'b0 | n3256_o;
  /* decoder.vhd:1434:13  */
  assign n3265_o = n3258_o ? 1'b1 : n2030_o;
  /* decoder.vhd:1434:13  */
  assign n3268_o = n3258_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1434:13  */
  assign n3271_o = n3258_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1433:11  */
  assign n3273_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1440:11  */
  assign n3275_o = clk_mstate_i == 3'b100;
  assign n3276_o = {n3275_o, n3273_o};
  /* decoder.vhd:1431:9  */
  always @*
    case (n3276_o)
      2'b10: n3279_o = 1'b1;
      2'b01: n3279_o = 1'b0;
      default: n3279_o = 1'b0;
    endcase
  /* decoder.vhd:1431:9  */
  always @*
    case (n3276_o)
      2'b10: n3280_o = n2030_o;
      2'b01: n3280_o = n3265_o;
      default: n3280_o = n2030_o;
    endcase
  /* decoder.vhd:1431:9  */
  always @*
    case (n3276_o)
      2'b10: n3282_o = 1'b0;
      2'b01: n3282_o = n3268_o;
      default: n3282_o = 1'b0;
    endcase
  /* decoder.vhd:1431:9  */
  always @*
    case (n3276_o)
      2'b10: n3284_o = 2'b01;
      2'b01: n3284_o = n3271_o;
      default: n3284_o = 2'b01;
    endcase
  /* decoder.vhd:1431:9  */
  always @*
    case (n3276_o)
      2'b10: n3287_o = 1'b1;
      2'b01: n3287_o = 1'b0;
      default: n3287_o = 1'b0;
    endcase
  /* decoder.vhd:1430:7  */
  assign n3289_o = opc_mnemonic_s == 6'b100011;
  /* decoder.vhd:1454:12  */
  assign n3290_o = ~clk_second_cycle_i;
  /* decoder.vhd:1454:52  */
  assign n3292_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1454:35  */
  assign n3293_o = n3292_o & n3290_o;
  /* decoder.vhd:1456:26  */
  assign n3294_o = opc_opcode_q[3];
  /* decoder.vhd:1456:30  */
  assign n3295_o = ~n3294_o;
  /* decoder.vhd:1455:42  */
  assign n3297_o = 1'b0 | n3295_o;
  /* decoder.vhd:1454:9  */
  assign n3304_o = n3311_o ? 1'b1 : n2030_o;
  /* decoder.vhd:1455:11  */
  assign n3307_o = n3297_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1455:11  */
  assign n3310_o = n3297_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1454:9  */
  assign n3311_o = n3293_o & n3297_o;
  /* decoder.vhd:1454:9  */
  assign n3313_o = n3293_o ? n3307_o : 1'b0;
  /* decoder.vhd:1454:9  */
  assign n3315_o = n3293_o ? n3310_o : 2'b01;
  /* decoder.vhd:1463:48  */
  assign n3317_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1463:31  */
  assign n3318_o = n3317_o & clk_second_cycle_i;
  /* decoder.vhd:1463:9  */
  assign n3321_o = n3318_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1450:7  */
  assign n3323_o = opc_mnemonic_s == 6'b100100;
  /* decoder.vhd:1470:25  */
  assign n3325_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1470:9  */
  assign n3328_o = n3325_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1470:9  */
  assign n3331_o = n3325_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1468:7  */
  assign n3333_o = opc_mnemonic_s == 6'b111111;
  /* decoder.vhd:1478:25  */
  assign n3335_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1479:26  */
  assign n3336_o = opc_opcode_q[5];
  /* decoder.vhd:1479:11  */
  assign n3339_o = n3336_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1479:11  */
  assign n3342_o = n3336_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1479:11  */
  assign n3345_o = n3336_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1479:11  */
  assign n3348_o = n3336_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1478:9  */
  assign n3350_o = n3335_o ? n3339_o : 1'b0;
  /* decoder.vhd:1478:9  */
  assign n3352_o = n3335_o ? n3342_o : 1'b0;
  /* decoder.vhd:1478:9  */
  assign n3354_o = n3335_o ? n3345_o : 1'b0;
  /* decoder.vhd:1478:9  */
  assign n3356_o = n3335_o ? n3348_o : 1'b0;
  /* decoder.vhd:1477:7  */
  assign n3358_o = opc_mnemonic_s == 6'b100101;
  /* decoder.vhd:1492:12  */
  assign n3359_o = ~clk_second_cycle_i;
  /* decoder.vhd:1498:53  */
  assign n3361_o = opc_opcode_q[1:0];
  /* decoder.vhd:1500:32  */
  assign n3362_o = opc_opcode_q[7:4];
  /* decoder.vhd:1501:17  */
  assign n3365_o = n3362_o == 4'b1001;
  /* decoder.vhd:1503:17  */
  assign n3368_o = n3362_o == 4'b1000;
  /* decoder.vhd:1505:17  */
  assign n3371_o = n3362_o == 4'b0011;
  assign n3372_o = {n3371_o, n3368_o, n3365_o};
  assign n3373_o = n2032_o[3:2];
  assign n3374_o = n2033_o[3:2];
  /* decoder.vhd:622:5  */
  assign n3375_o = n2019_o ? n3373_o : n3374_o;
  /* decoder.vhd:1500:15  */
  always @*
    case (n3372_o)
      3'b100: n3376_o = 2'b01;
      3'b010: n3376_o = 2'b10;
      3'b001: n3376_o = 2'b11;
      default: n3376_o = n3375_o;
    endcase
  /* decoder.vhd:1495:13  */
  assign n3378_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1516:13  */
  assign n3380_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1522:13  */
  assign n3382_o = clk_mstate_i == 3'b100;
  assign n3383_o = {n3382_o, n3380_o, n3378_o};
  /* decoder.vhd:1493:11  */
  always @*
    case (n3383_o)
      3'b100: n3386_o = 1'b0;
      3'b010: n3386_o = 1'b1;
      3'b001: n3386_o = 1'b0;
      default: n3386_o = 1'b0;
    endcase
  /* decoder.vhd:1493:11  */
  always @*
    case (n3383_o)
      3'b100: n3390_o = 1'b0;
      3'b010: n3390_o = 1'b1;
      3'b001: n3390_o = 1'b1;
      default: n3390_o = 1'b0;
    endcase
  assign n3391_o = n2032_o[1:0];
  assign n3392_o = n2033_o[1:0];
  /* decoder.vhd:622:5  */
  assign n3393_o = n2019_o ? n3391_o : n3392_o;
  /* decoder.vhd:1493:11  */
  always @*
    case (n3383_o)
      3'b100: n3394_o = n3393_o;
      3'b010: n3394_o = n3393_o;
      3'b001: n3394_o = n3361_o;
      default: n3394_o = n3393_o;
    endcase
  assign n3395_o = n2032_o[3:2];
  assign n3396_o = n2033_o[3:2];
  /* decoder.vhd:622:5  */
  assign n3397_o = n2019_o ? n3395_o : n3396_o;
  /* decoder.vhd:1493:11  */
  always @*
    case (n3383_o)
      3'b100: n3398_o = n3397_o;
      3'b010: n3398_o = n3397_o;
      3'b001: n3398_o = n3376_o;
      default: n3398_o = n3397_o;
    endcase
  assign n3399_o = n2032_o[7:4];
  assign n3400_o = n2033_o[7:4];
  /* decoder.vhd:622:5  */
  assign n3401_o = n2019_o ? n3399_o : n3400_o;
  /* decoder.vhd:1493:11  */
  always @*
    case (n3383_o)
      3'b100: n3402_o = n3401_o;
      3'b010: n3402_o = n3401_o;
      3'b001: n3402_o = 4'b0000;
      default: n3402_o = n3401_o;
    endcase
  /* decoder.vhd:1493:11  */
  always @*
    case (n3383_o)
      3'b100: n3404_o = n2038_o;
      3'b010: n3404_o = n2038_o;
      3'b001: n3404_o = 1'b1;
      default: n3404_o = n2038_o;
    endcase
  /* decoder.vhd:1493:11  */
  always @*
    case (n3383_o)
      3'b100: n3408_o = 1'b1;
      3'b010: n3408_o = 1'b1;
      3'b001: n3408_o = 1'b0;
      default: n3408_o = 1'b0;
    endcase
  /* decoder.vhd:1532:27  */
  assign n3410_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1532:53  */
  assign n3412_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1532:37  */
  assign n3413_o = n3410_o | n3412_o;
  /* decoder.vhd:1532:11  */
  assign n3416_o = n3413_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1492:9  */
  assign n3418_o = n3359_o ? n3386_o : 1'b0;
  /* decoder.vhd:1492:9  */
  assign n3420_o = n3359_o ? n3390_o : 1'b0;
  assign n3421_o = {n3402_o, n3398_o, n3394_o};
  /* decoder.vhd:1492:9  */
  assign n3422_o = n3359_o ? n3421_o : n2034_o;
  /* decoder.vhd:1492:9  */
  assign n3423_o = n3359_o ? n3404_o : n2038_o;
  /* decoder.vhd:1492:9  */
  assign n3424_o = n3359_o ? n3408_o : n3416_o;
  /* decoder.vhd:1489:7  */
  assign n3426_o = opc_mnemonic_s == 6'b101101;
  /* decoder.vhd:1542:12  */
  assign n3427_o = ~clk_second_cycle_i;
  /* decoder.vhd:1548:53  */
  assign n3428_o = opc_opcode_q[1:0];
  /* decoder.vhd:1547:48  */
  assign n3430_o = {6'b000000, n3428_o};
  /* decoder.vhd:1545:13  */
  assign n3432_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1554:13  */
  assign n3435_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1561:13  */
  assign n3437_o = clk_mstate_i == 3'b100;
  assign n3438_o = {n3437_o, n3435_o, n3432_o};
  /* decoder.vhd:1543:11  */
  always @*
    case (n3438_o)
      3'b100: n3442_o = 1'b0;
      3'b010: n3442_o = 1'b1;
      3'b001: n3442_o = 1'b1;
      default: n3442_o = 1'b0;
    endcase
  assign n3443_o = n3430_o[3:0];
  assign n3444_o = n2032_o[3:0];
  assign n3445_o = n2033_o[3:0];
  /* decoder.vhd:622:5  */
  assign n3446_o = n2019_o ? n3444_o : n3445_o;
  /* decoder.vhd:1543:11  */
  always @*
    case (n3438_o)
      3'b100: n3447_o = n3446_o;
      3'b010: n3447_o = 4'b1111;
      3'b001: n3447_o = n3443_o;
      default: n3447_o = n3446_o;
    endcase
  assign n3448_o = n3430_o[7:4];
  assign n3449_o = n2032_o[7:4];
  assign n3450_o = n2033_o[7:4];
  /* decoder.vhd:622:5  */
  assign n3451_o = n2019_o ? n3449_o : n3450_o;
  /* decoder.vhd:1543:11  */
  always @*
    case (n3438_o)
      3'b100: n3452_o = n3451_o;
      3'b010: n3452_o = n3451_o;
      3'b001: n3452_o = n3448_o;
      default: n3452_o = n3451_o;
    endcase
  /* decoder.vhd:1543:11  */
  always @*
    case (n3438_o)
      3'b100: n3455_o = n2038_o;
      3'b010: n3455_o = 1'b1;
      3'b001: n3455_o = 1'b1;
      default: n3455_o = n2038_o;
    endcase
  /* decoder.vhd:1543:11  */
  always @*
    case (n3438_o)
      3'b100: n3459_o = 1'b1;
      3'b010: n3459_o = 1'b1;
      3'b001: n3459_o = 1'b0;
      default: n3459_o = 1'b0;
    endcase
  /* decoder.vhd:1572:13  */
  assign n3461_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1577:13  */
  assign n3463_o = clk_mstate_i == 3'b001;
  assign n3464_o = {n3463_o, n3461_o};
  /* decoder.vhd:1570:11  */
  always @*
    case (n3464_o)
      2'b10: n3467_o = 1'b1;
      2'b01: n3467_o = 1'b0;
      default: n3467_o = 1'b0;
    endcase
  /* decoder.vhd:1570:11  */
  always @*
    case (n3464_o)
      2'b10: n3470_o = 1'b1;
      2'b01: n3470_o = 1'b0;
      default: n3470_o = 1'b0;
    endcase
  /* decoder.vhd:1570:11  */
  always @*
    case (n3464_o)
      2'b10: n3473_o = 1'b1;
      2'b01: n3473_o = 1'b0;
      default: n3473_o = 1'b0;
    endcase
  /* decoder.vhd:1570:11  */
  always @*
    case (n3464_o)
      2'b10: n3477_o = 1'b1;
      2'b01: n3477_o = 1'b1;
      default: n3477_o = 1'b0;
    endcase
  /* decoder.vhd:1542:9  */
  assign n3479_o = n3427_o ? 1'b0 : n3467_o;
  /* decoder.vhd:1542:9  */
  assign n3481_o = n3427_o ? n3442_o : 1'b0;
  /* decoder.vhd:1542:9  */
  assign n3483_o = n3427_o ? 1'b0 : n3470_o;
  /* decoder.vhd:1542:9  */
  assign n3485_o = n3427_o ? 1'b0 : n3473_o;
  assign n3486_o = {n3452_o, n3447_o};
  /* decoder.vhd:1542:9  */
  assign n3487_o = n3427_o ? n3486_o : n2034_o;
  /* decoder.vhd:1542:9  */
  assign n3488_o = n3427_o ? n3455_o : n2038_o;
  /* decoder.vhd:1542:9  */
  assign n3489_o = n3427_o ? n3459_o : n3477_o;
  /* decoder.vhd:1539:7  */
  assign n3491_o = opc_mnemonic_s == 6'b100110;
  /* decoder.vhd:1594:12  */
  assign n3492_o = ~clk_second_cycle_i;
  /* decoder.vhd:1597:27  */
  assign n3494_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1599:28  */
  assign n3495_o = opc_opcode_q[6];
  /* decoder.vhd:1599:32  */
  assign n3496_o = ~n3495_o;
  /* decoder.vhd:1599:13  */
  assign n3499_o = n3496_o ? 2'b01 : 2'b10;
  /* decoder.vhd:1597:11  */
  assign n3502_o = n3494_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1597:11  */
  assign n3504_o = n3494_o ? n3499_o : 2'b00;
  /* decoder.vhd:1607:27  */
  assign n3506_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1607:11  */
  assign n3509_o = n3506_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1607:11  */
  assign n3512_o = n3506_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1594:9  */
  assign n3514_o = n3492_o ? 1'b0 : n3509_o;
  /* decoder.vhd:1594:9  */
  assign n3516_o = n3492_o ? n3502_o : 1'b0;
  /* decoder.vhd:1594:9  */
  assign n3518_o = n3492_o ? n3504_o : 2'b00;
  /* decoder.vhd:1594:9  */
  assign n3520_o = n3492_o ? 1'b0 : n3512_o;
  /* decoder.vhd:1591:7  */
  assign n3522_o = opc_mnemonic_s == 6'b100111;
  /* decoder.vhd:1621:24  */
  assign n3523_o = opc_opcode_q[4];
  /* decoder.vhd:1621:28  */
  assign n3524_o = ~n3523_o;
  /* decoder.vhd:1621:9  */
  assign n3527_o = n3524_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1621:9  */
  assign n3530_o = n3524_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1627:12  */
  assign n3531_o = ~clk_second_cycle_i;
  /* decoder.vhd:1631:13  */
  assign n3533_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1637:30  */
  assign n3534_o = opc_opcode_q[4];
  /* decoder.vhd:1637:15  */
  assign n3537_o = n3534_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1637:15  */
  assign n3540_o = n3534_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1636:13  */
  assign n3542_o = clk_mstate_i == 3'b100;
  assign n3543_o = {n3542_o, n3533_o};
  /* decoder.vhd:1629:11  */
  always @*
    case (n3543_o)
      2'b10: n3545_o = n3537_o;
      2'b01: n3545_o = 1'b0;
      default: n3545_o = 1'b0;
    endcase
  /* decoder.vhd:1629:11  */
  always @*
    case (n3543_o)
      2'b10: n3548_o = n3540_o;
      2'b01: n3548_o = 1'b1;
      default: n3548_o = 1'b0;
    endcase
  /* decoder.vhd:1629:11  */
  always @*
    case (n3543_o)
      2'b10: n3551_o = 1'b0;
      2'b01: n3551_o = 1'b1;
      default: n3551_o = 1'b0;
    endcase
  /* decoder.vhd:1647:27  */
  assign n3553_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1648:28  */
  assign n3554_o = opc_opcode_q[4];
  /* decoder.vhd:1648:32  */
  assign n3555_o = ~n3554_o;
  /* decoder.vhd:1648:13  */
  assign n3558_o = n3555_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1648:13  */
  assign n3561_o = n3555_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1648:13  */
  assign n3564_o = n3555_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1648:13  */
  assign n3567_o = n3555_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1647:11  */
  assign n3569_o = n3553_o ? n3558_o : 1'b0;
  /* decoder.vhd:1647:11  */
  assign n3571_o = n3553_o ? n3561_o : 1'b0;
  /* decoder.vhd:1647:11  */
  assign n3573_o = n3553_o ? n3564_o : 1'b0;
  /* decoder.vhd:1647:11  */
  assign n3575_o = n3553_o ? n3567_o : 1'b0;
  /* decoder.vhd:1627:9  */
  assign n3577_o = n3531_o ? 1'b0 : n3569_o;
  /* decoder.vhd:1627:9  */
  assign n3578_o = n3531_o ? n3545_o : n3571_o;
  /* decoder.vhd:1627:9  */
  assign n3579_o = n3531_o ? n3548_o : n3573_o;
  /* decoder.vhd:1627:9  */
  assign n3581_o = n3531_o ? n3551_o : 1'b0;
  /* decoder.vhd:1627:9  */
  assign n3583_o = n3531_o ? 1'b0 : n3575_o;
  /* decoder.vhd:1627:9  */
  assign n3586_o = n3531_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1618:7  */
  assign n3588_o = opc_mnemonic_s == 6'b101000;
  /* decoder.vhd:1663:7  */
  assign n3590_o = opc_mnemonic_s == 6'b101001;
  /* decoder.vhd:1672:28  */
  assign n3591_o = opc_opcode_q[3];
  /* decoder.vhd:1672:32  */
  assign n3592_o = ~n3591_o;
  /* decoder.vhd:1671:44  */
  assign n3594_o = 1'b0 | n3592_o;
  /* decoder.vhd:1671:13  */
  assign n3601_o = n3594_o ? 1'b1 : n2030_o;
  /* decoder.vhd:1671:13  */
  assign n3604_o = n3594_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1671:13  */
  assign n3607_o = n3594_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1670:11  */
  assign n3609_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1677:11  */
  assign n3614_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1681:11  */
  assign n3619_o = clk_mstate_i == 3'b100;
  assign n3620_o = {n3619_o, n3614_o, n3609_o};
  /* decoder.vhd:1668:9  */
  always @*
    case (n3620_o)
      3'b100: n3623_o = 1'b1;
      3'b010: n3623_o = 1'b0;
      3'b001: n3623_o = 1'b0;
      default: n3623_o = 1'b0;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3620_o)
      3'b100: n3626_o = 1'b0;
      3'b010: n3626_o = 1'b1;
      3'b001: n3626_o = 1'b0;
      default: n3626_o = 1'b0;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3620_o)
      3'b100: n3629_o = 1'b1;
      3'b010: n3629_o = 1'b0;
      3'b001: n3629_o = 1'b0;
      default: n3629_o = 1'b0;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3620_o)
      3'b100: n3630_o = n2030_o;
      3'b010: n3630_o = n2030_o;
      3'b001: n3630_o = n3601_o;
      default: n3630_o = n2030_o;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3620_o)
      3'b100: n3633_o = 1'b0;
      3'b010: n3633_o = 1'b1;
      3'b001: n3633_o = n3604_o;
      default: n3633_o = 1'b0;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3620_o)
      3'b100: n3636_o = 4'b0001;
      3'b010: n3636_o = 4'b1100;
      3'b001: n3636_o = 4'b1100;
      default: n3636_o = 4'b1100;
    endcase
  /* decoder.vhd:1668:9  */
  always @*
    case (n3620_o)
      3'b100: n3638_o = 2'b01;
      3'b010: n3638_o = 2'b01;
      3'b001: n3638_o = n3607_o;
      default: n3638_o = 2'b01;
    endcase
  /* decoder.vhd:1667:7  */
  assign n3640_o = opc_mnemonic_s == 6'b101010;
  /* decoder.vhd:1696:13  */
  assign n3642_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1700:13  */
  assign n3647_o = clk_mstate_i == 3'b010;
  assign n3648_o = {n3647_o, n3642_o};
  /* decoder.vhd:1694:11  */
  always @*
    case (n3648_o)
      2'b10: n3651_o = 1'b1;
      2'b01: n3651_o = 1'b0;
      default: n3651_o = 1'b0;
    endcase
  /* decoder.vhd:1694:11  */
  always @*
    case (n3648_o)
      2'b10: n3654_o = 1'b0;
      2'b01: n3654_o = 1'b1;
      default: n3654_o = 1'b0;
    endcase
  /* decoder.vhd:1694:11  */
  always @*
    case (n3648_o)
      2'b10: n3657_o = 1'b1;
      2'b01: n3657_o = 1'b0;
      default: n3657_o = 1'b0;
    endcase
  /* decoder.vhd:1694:11  */
  always @*
    case (n3648_o)
      2'b10: n3660_o = 4'b0001;
      2'b01: n3660_o = 4'b1100;
      default: n3660_o = 4'b1100;
    endcase
  /* decoder.vhd:1693:9  */
  assign n3662_o = clk_second_cycle_i ? n3651_o : 1'b0;
  /* decoder.vhd:1693:9  */
  assign n3664_o = clk_second_cycle_i ? n3654_o : 1'b0;
  /* decoder.vhd:1693:9  */
  assign n3666_o = clk_second_cycle_i ? n3657_o : 1'b0;
  /* decoder.vhd:1693:9  */
  assign n3668_o = clk_second_cycle_i ? n3660_o : 4'b1100;
  /* decoder.vhd:1690:7  */
  assign n3670_o = opc_mnemonic_s == 6'b101011;
  /* decoder.vhd:1714:12  */
  assign n3671_o = ~clk_second_cycle_i;
  /* decoder.vhd:1716:27  */
  assign n3673_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:1717:28  */
  assign n3674_o = opc_opcode_q[1:0];
  /* decoder.vhd:1717:41  */
  assign n3676_o = n3674_o == 2'b00;
  /* decoder.vhd:1719:31  */
  assign n3677_o = opc_opcode_q[1];
  /* decoder.vhd:1719:35  */
  assign n3678_o = ~n3677_o;
  /* decoder.vhd:1719:13  */
  assign n3681_o = n3678_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1719:13  */
  assign n3684_o = n3678_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1719:13  */
  assign n3687_o = n3678_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1719:13  */
  assign n3690_o = n3678_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1717:13  */
  assign n3692_o = n3676_o ? 1'b0 : n3681_o;
  /* decoder.vhd:1717:13  */
  assign n3694_o = n3676_o ? 1'b0 : n3684_o;
  /* decoder.vhd:1717:13  */
  assign n3696_o = n3676_o ? 1'b0 : n3687_o;
  /* decoder.vhd:1717:13  */
  assign n3698_o = n3676_o ? 1'b0 : n3690_o;
  /* decoder.vhd:1717:13  */
  assign n3701_o = n3676_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3704_o = n3673_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3706_o = n3673_o ? n3692_o : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3708_o = n3673_o ? n3694_o : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3710_o = n3673_o ? n3696_o : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3712_o = n3673_o ? n3698_o : 1'b0;
  /* decoder.vhd:1716:11  */
  assign n3714_o = n3673_o ? n3701_o : 1'b0;
  /* decoder.vhd:1734:13  */
  assign n3716_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1739:13  */
  assign n3718_o = clk_mstate_i == 3'b001;
  /* decoder.vhd:1748:30  */
  assign n3719_o = opc_opcode_q[1:0];
  /* decoder.vhd:1748:43  */
  assign n3721_o = n3719_o == 2'b00;
  /* decoder.vhd:1750:33  */
  assign n3722_o = opc_opcode_q[1];
  /* decoder.vhd:1750:37  */
  assign n3723_o = ~n3722_o;
  /* decoder.vhd:1750:15  */
  assign n3726_o = n3723_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1750:15  */
  assign n3729_o = n3723_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1748:15  */
  assign n3732_o = n3721_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1748:15  */
  assign n3734_o = n3721_o ? 1'b0 : n3726_o;
  /* decoder.vhd:1748:15  */
  assign n3736_o = n3721_o ? 1'b0 : n3729_o;
  /* decoder.vhd:1744:13  */
  assign n3738_o = clk_mstate_i == 3'b010;
  assign n3739_o = {n3738_o, n3718_o, n3716_o};
  /* decoder.vhd:1731:11  */
  always @*
    case (n3739_o)
      3'b100: n3743_o = 1'b0;
      3'b010: n3743_o = 1'b1;
      3'b001: n3743_o = 1'b1;
      default: n3743_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3739_o)
      3'b100: n3747_o = 1'b1;
      3'b010: n3747_o = 1'b1;
      3'b001: n3747_o = 1'b0;
      default: n3747_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3739_o)
      3'b100: n3749_o = n3732_o;
      3'b010: n3749_o = 1'b0;
      3'b001: n3749_o = 1'b0;
      default: n3749_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3739_o)
      3'b100: n3751_o = n3734_o;
      3'b010: n3751_o = 1'b0;
      3'b001: n3751_o = 1'b0;
      default: n3751_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3739_o)
      3'b100: n3753_o = n3736_o;
      3'b010: n3753_o = 1'b0;
      3'b001: n3753_o = 1'b0;
      default: n3753_o = 1'b0;
    endcase
  /* decoder.vhd:1731:11  */
  always @*
    case (n3739_o)
      3'b100: n3756_o = 4'b0001;
      3'b010: n3756_o = 4'b1100;
      3'b001: n3756_o = 4'b1100;
      default: n3756_o = 4'b1100;
    endcase
  /* decoder.vhd:1714:9  */
  assign n3758_o = n3671_o ? 1'b0 : n3743_o;
  /* decoder.vhd:1714:9  */
  assign n3760_o = n3671_o ? n3704_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3762_o = n3671_o ? 1'b0 : n3747_o;
  /* decoder.vhd:1714:9  */
  assign n3764_o = n3671_o ? 1'b0 : n3749_o;
  /* decoder.vhd:1714:9  */
  assign n3766_o = n3671_o ? 1'b0 : n3751_o;
  /* decoder.vhd:1714:9  */
  assign n3768_o = n3671_o ? n3706_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3770_o = n3671_o ? 1'b0 : n3753_o;
  /* decoder.vhd:1714:9  */
  assign n3772_o = n3671_o ? n3708_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3774_o = n3671_o ? 4'b1100 : n3756_o;
  /* decoder.vhd:1714:9  */
  assign n3776_o = n3671_o ? n3710_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3778_o = n3671_o ? n3712_o : 1'b0;
  /* decoder.vhd:1714:9  */
  assign n3780_o = n3671_o ? n3714_o : 1'b0;
  /* decoder.vhd:1711:7  */
  assign n3782_o = opc_mnemonic_s == 6'b101100;
  /* decoder.vhd:1766:25  */
  assign n3784_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1766:9  */
  assign n3787_o = n3784_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1766:9  */
  assign n3790_o = n3784_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1764:7  */
  assign n3792_o = opc_mnemonic_s == 6'b111011;
  /* decoder.vhd:1774:24  */
  assign n3793_o = opc_opcode_q[4];
  /* decoder.vhd:1774:28  */
  assign n3794_o = ~n3793_o;
  /* decoder.vhd:1774:9  */
  assign n3797_o = n3794_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1779:12  */
  assign n3798_o = ~clk_second_cycle_i;
  /* decoder.vhd:1779:52  */
  assign n3800_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1779:35  */
  assign n3801_o = n3800_o & n3798_o;
  /* decoder.vhd:1782:26  */
  assign n3802_o = opc_opcode_q[4];
  /* decoder.vhd:1783:28  */
  assign n3803_o = opc_opcode_q[1];
  /* decoder.vhd:1783:32  */
  assign n3804_o = ~n3803_o;
  /* decoder.vhd:1783:13  */
  assign n3807_o = n3804_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1783:13  */
  assign n3810_o = n3804_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1782:11  */
  assign n3813_o = n3802_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1782:11  */
  assign n3815_o = n3802_o ? n3807_o : 1'b0;
  /* decoder.vhd:1782:11  */
  assign n3817_o = n3802_o ? n3810_o : 1'b0;
  /* decoder.vhd:1779:9  */
  assign n3820_o = n3801_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1779:9  */
  assign n3822_o = n3801_o ? n3813_o : 1'b0;
  /* decoder.vhd:1779:9  */
  assign n3824_o = n3801_o ? n3815_o : 1'b0;
  /* decoder.vhd:1779:9  */
  assign n3826_o = n3801_o ? n3817_o : 1'b0;
  /* decoder.vhd:1773:7  */
  assign n3828_o = opc_mnemonic_s == 6'b101110;
  /* decoder.vhd:1798:12  */
  assign n3829_o = ~clk_second_cycle_i;
  /* decoder.vhd:1801:13  */
  assign n3831_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1805:13  */
  assign n3833_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1812:13  */
  assign n3835_o = clk_mstate_i == 3'b100;
  assign n3836_o = {n3835_o, n3833_o, n3831_o};
  /* decoder.vhd:1799:11  */
  always @*
    case (n3836_o)
      3'b100: n3839_o = 1'b1;
      3'b010: n3839_o = 1'b1;
      3'b001: n3839_o = n2030_o;
      default: n3839_o = n2030_o;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3836_o)
      3'b100: n3842_o = 1'b1;
      3'b010: n3842_o = 1'b0;
      3'b001: n3842_o = 1'b0;
      default: n3842_o = 1'b0;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3836_o)
      3'b100: n3845_o = 1'b1;
      3'b010: n3845_o = 1'b0;
      3'b001: n3845_o = 1'b0;
      default: n3845_o = 1'b0;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3836_o)
      3'b100: n3848_o = 1'b0;
      3'b010: n3848_o = 1'b1;
      3'b001: n3848_o = 1'b0;
      default: n3848_o = 1'b0;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3836_o)
      3'b100: n3852_o = 2'b11;
      3'b010: n3852_o = 2'b10;
      3'b001: n3852_o = 2'b01;
      default: n3852_o = 2'b01;
    endcase
  /* decoder.vhd:1799:11  */
  always @*
    case (n3836_o)
      3'b100: n3855_o = 1'b0;
      3'b010: n3855_o = 1'b0;
      3'b001: n3855_o = 1'b1;
      default: n3855_o = 1'b0;
    endcase
  /* decoder.vhd:1829:30  */
  assign n3856_o = opc_opcode_q[4];
  /* decoder.vhd:1829:15  */
  assign n3859_o = n3856_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1829:15  */
  assign n3862_o = n3856_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1826:13  */
  assign n3864_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1834:13  */
  assign n3866_o = clk_mstate_i == 3'b001;
  assign n3867_o = {n3866_o, n3864_o};
  /* decoder.vhd:1824:11  */
  always @*
    case (n3867_o)
      2'b10: n3870_o = 1'b0;
      2'b01: n3870_o = 1'b1;
      default: n3870_o = 1'b0;
    endcase
  /* decoder.vhd:1824:11  */
  always @*
    case (n3867_o)
      2'b10: n3873_o = 1'b0;
      2'b01: n3873_o = 1'b1;
      default: n3873_o = 1'b0;
    endcase
  /* decoder.vhd:1824:11  */
  always @*
    case (n3867_o)
      2'b10: n3875_o = 1'b0;
      2'b01: n3875_o = n3859_o;
      default: n3875_o = 1'b0;
    endcase
  /* decoder.vhd:1824:11  */
  always @*
    case (n3867_o)
      2'b10: n3878_o = 1'b1;
      2'b01: n3878_o = 1'b0;
      default: n3878_o = 1'b0;
    endcase
  /* decoder.vhd:1824:11  */
  always @*
    case (n3867_o)
      2'b10: n3880_o = 1'b0;
      2'b01: n3880_o = n3862_o;
      default: n3880_o = 1'b0;
    endcase
  /* decoder.vhd:1798:9  */
  assign n3881_o = n3829_o ? n3839_o : n2030_o;
  /* decoder.vhd:1798:9  */
  assign n3882_o = n3829_o ? n3842_o : n3870_o;
  /* decoder.vhd:1798:9  */
  assign n3884_o = n3829_o ? n3845_o : 1'b0;
  /* decoder.vhd:1798:9  */
  assign n3886_o = n3829_o ? 1'b0 : n3873_o;
  /* decoder.vhd:1798:9  */
  assign n3888_o = n3829_o ? n3848_o : 1'b0;
  /* decoder.vhd:1798:9  */
  assign n3890_o = n3829_o ? 1'b0 : n3875_o;
  /* decoder.vhd:1798:9  */
  assign n3892_o = n3829_o ? n3852_o : 2'b01;
  /* decoder.vhd:1798:9  */
  assign n3894_o = n3829_o ? n3855_o : 1'b0;
  /* decoder.vhd:1798:9  */
  assign n3896_o = n3829_o ? 1'b0 : n3878_o;
  /* decoder.vhd:1798:9  */
  assign n3898_o = n3829_o ? 1'b0 : n3880_o;
  /* decoder.vhd:1797:7  */
  assign n3900_o = opc_mnemonic_s == 6'b101111;
  /* decoder.vhd:1846:25  */
  assign n3902_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1851:26  */
  assign n3903_o = opc_opcode_q[4];
  /* decoder.vhd:1851:11  */
  assign n3906_o = n3903_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1851:11  */
  assign n3908_o = n3903_o ? alu_carry_i : 1'b0;
  /* decoder.vhd:1851:11  */
  assign n3911_o = n3903_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n3914_o = n3902_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n3917_o = n3902_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n3920_o = n3902_o ? 4'b0101 : 4'b1100;
  /* decoder.vhd:1846:9  */
  assign n3922_o = n3902_o ? n3906_o : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n3924_o = n3902_o ? n3908_o : 1'b0;
  /* decoder.vhd:1846:9  */
  assign n3926_o = n3902_o ? n3911_o : 1'b0;
  /* decoder.vhd:1845:7  */
  assign n3928_o = opc_mnemonic_s == 6'b110000;
  /* decoder.vhd:1860:25  */
  assign n3930_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1865:26  */
  assign n3931_o = opc_opcode_q[4];
  /* decoder.vhd:1865:30  */
  assign n3932_o = ~n3931_o;
  /* decoder.vhd:1865:11  */
  assign n3935_o = n3932_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1865:11  */
  assign n3937_o = n3932_o ? alu_carry_i : 1'b0;
  /* decoder.vhd:1865:11  */
  assign n3940_o = n3932_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n3943_o = n3930_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n3946_o = n3930_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n3949_o = n3930_o ? 4'b0110 : 4'b1100;
  /* decoder.vhd:1860:9  */
  assign n3951_o = n3930_o ? n3935_o : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n3953_o = n3930_o ? n3937_o : 1'b0;
  /* decoder.vhd:1860:9  */
  assign n3955_o = n3930_o ? n3940_o : 1'b0;
  /* decoder.vhd:1859:7  */
  assign n3957_o = opc_mnemonic_s == 6'b110001;
  /* decoder.vhd:1874:25  */
  assign n3959_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1875:26  */
  assign n3960_o = opc_opcode_q[4];
  /* decoder.vhd:1875:11  */
  assign n3963_o = n3960_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1875:11  */
  assign n3966_o = n3960_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1874:9  */
  assign n3968_o = n3959_o ? n3963_o : 1'b0;
  /* decoder.vhd:1874:9  */
  assign n3970_o = n3959_o ? n3966_o : 1'b0;
  /* decoder.vhd:1873:7  */
  assign n3972_o = opc_mnemonic_s == 6'b110010;
  /* decoder.vhd:1884:25  */
  assign n3974_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1885:45  */
  assign n3975_o = opc_opcode_q[4];
  /* decoder.vhd:1884:9  */
  assign n3977_o = n3974_o ? n3975_o : 1'b0;
  /* decoder.vhd:1884:9  */
  assign n3980_o = n3974_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1883:7  */
  assign n3982_o = opc_mnemonic_s == 6'b110011;
  /* decoder.vhd:1891:25  */
  assign n3984_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1891:9  */
  assign n3987_o = n3984_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1890:7  */
  assign n3989_o = opc_mnemonic_s == 6'b110100;
  /* decoder.vhd:1897:25  */
  assign n3991_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1898:26  */
  assign n3992_o = opc_opcode_q[4];
  /* decoder.vhd:1898:11  */
  assign n3995_o = n3992_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1898:11  */
  assign n3998_o = n3992_o ? 1'b0 : 1'b1;
  /* decoder.vhd:1897:9  */
  assign n4000_o = n3991_o ? n3995_o : 1'b0;
  /* decoder.vhd:1897:9  */
  assign n4002_o = n3991_o ? n3998_o : 1'b0;
  /* decoder.vhd:1896:7  */
  assign n4004_o = opc_mnemonic_s == 6'b110101;
  /* decoder.vhd:1909:25  */
  assign n4006_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1909:9  */
  assign n4009_o = n4006_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1909:9  */
  assign n4012_o = n4006_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1906:7  */
  assign n4014_o = opc_mnemonic_s == 6'b110110;
  /* decoder.vhd:1920:28  */
  assign n4015_o = opc_opcode_q[3];
  /* decoder.vhd:1920:32  */
  assign n4016_o = ~n4015_o;
  /* decoder.vhd:1919:44  */
  assign n4018_o = 1'b0 | n4016_o;
  /* decoder.vhd:1919:13  */
  assign n4025_o = n4018_o ? 1'b1 : n2030_o;
  /* decoder.vhd:1919:13  */
  assign n4028_o = n4018_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1919:13  */
  assign n4031_o = n4018_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1918:11  */
  assign n4033_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1930:28  */
  assign n4034_o = opc_opcode_q[4];
  /* decoder.vhd:1930:13  */
  assign n4037_o = n4034_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1926:11  */
  assign n4039_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1940:28  */
  assign n4040_o = opc_opcode_q[4];
  /* decoder.vhd:1940:13  */
  assign n4043_o = n4040_o ? 4'b1011 : 4'b1100;
  /* decoder.vhd:1937:11  */
  assign n4045_o = clk_mstate_i == 3'b100;
  assign n4046_o = {n4045_o, n4039_o, n4033_o};
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4049_o = 1'b0;
      3'b010: n4049_o = 1'b1;
      3'b001: n4049_o = 1'b0;
      default: n4049_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4052_o = 1'b0;
      3'b010: n4052_o = 1'b1;
      3'b001: n4052_o = 1'b0;
      default: n4052_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4055_o = 1'b1;
      3'b010: n4055_o = 1'b0;
      3'b001: n4055_o = 1'b0;
      default: n4055_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4056_o = n2030_o;
      3'b010: n4056_o = n2030_o;
      3'b001: n4056_o = n4025_o;
      default: n4056_o = n2030_o;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4059_o = 1'b0;
      3'b010: n4059_o = 1'b1;
      3'b001: n4059_o = n4028_o;
      default: n4059_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4061_o = n4043_o;
      3'b010: n4061_o = 4'b1100;
      3'b001: n4061_o = 4'b1100;
      default: n4061_o = 4'b1100;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4063_o = 1'b0;
      3'b010: n4063_o = n4037_o;
      3'b001: n4063_o = 1'b0;
      default: n4063_o = 1'b0;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4065_o = 2'b01;
      3'b010: n4065_o = 2'b01;
      3'b001: n4065_o = n4031_o;
      default: n4065_o = 2'b01;
    endcase
  /* decoder.vhd:1916:9  */
  always @*
    case (n4046_o)
      3'b100: n4068_o = 1'b1;
      3'b010: n4068_o = 1'b0;
      3'b001: n4068_o = 1'b0;
      default: n4068_o = 1'b0;
    endcase
  /* decoder.vhd:1915:7  */
  assign n4070_o = opc_mnemonic_s == 6'b110111;
  /* decoder.vhd:1957:28  */
  assign n4071_o = opc_opcode_q[3];
  /* decoder.vhd:1957:32  */
  assign n4072_o = ~n4071_o;
  /* decoder.vhd:1956:44  */
  assign n4074_o = 1'b0 | n4072_o;
  /* decoder.vhd:1956:13  */
  assign n4081_o = n4074_o ? 1'b1 : n2030_o;
  /* decoder.vhd:1956:13  */
  assign n4084_o = n4074_o ? 1'b1 : 1'b0;
  /* decoder.vhd:1956:13  */
  assign n4087_o = n4074_o ? 2'b00 : 2'b01;
  /* decoder.vhd:1955:11  */
  assign n4089_o = clk_mstate_i == 3'b010;
  /* decoder.vhd:1962:11  */
  assign n4094_o = clk_mstate_i == 3'b011;
  /* decoder.vhd:1966:11  */
  assign n4099_o = clk_mstate_i == 3'b100;
  assign n4100_o = {n4099_o, n4094_o, n4089_o};
  /* decoder.vhd:1953:9  */
  always @*
    case (n4100_o)
      3'b100: n4103_o = 1'b1;
      3'b010: n4103_o = 1'b0;
      3'b001: n4103_o = 1'b0;
      default: n4103_o = 1'b0;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4100_o)
      3'b100: n4106_o = 1'b0;
      3'b010: n4106_o = 1'b1;
      3'b001: n4106_o = 1'b0;
      default: n4106_o = 1'b0;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4100_o)
      3'b100: n4109_o = 1'b1;
      3'b010: n4109_o = 1'b0;
      3'b001: n4109_o = 1'b0;
      default: n4109_o = 1'b0;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4100_o)
      3'b100: n4110_o = n2030_o;
      3'b010: n4110_o = n2030_o;
      3'b001: n4110_o = n4081_o;
      default: n4110_o = n2030_o;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4100_o)
      3'b100: n4113_o = 1'b0;
      3'b010: n4113_o = 1'b1;
      3'b001: n4113_o = n4084_o;
      default: n4113_o = 1'b0;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4100_o)
      3'b100: n4116_o = 4'b0010;
      3'b010: n4116_o = 4'b1100;
      3'b001: n4116_o = 4'b1100;
      default: n4116_o = 4'b1100;
    endcase
  /* decoder.vhd:1953:9  */
  always @*
    case (n4100_o)
      3'b100: n4118_o = 2'b01;
      3'b010: n4118_o = 2'b01;
      3'b001: n4118_o = n4087_o;
      default: n4118_o = 2'b01;
    endcase
  /* decoder.vhd:1952:7  */
  assign n4120_o = opc_mnemonic_s == 6'b111000;
  /* decoder.vhd:1981:13  */
  assign n4122_o = clk_mstate_i == 3'b000;
  /* decoder.vhd:1985:13  */
  assign n4127_o = clk_mstate_i == 3'b010;
  assign n4128_o = {n4127_o, n4122_o};
  /* decoder.vhd:1979:11  */
  always @*
    case (n4128_o)
      2'b10: n4131_o = 1'b1;
      2'b01: n4131_o = 1'b0;
      default: n4131_o = 1'b0;
    endcase
  /* decoder.vhd:1979:11  */
  always @*
    case (n4128_o)
      2'b10: n4134_o = 1'b0;
      2'b01: n4134_o = 1'b1;
      default: n4134_o = 1'b0;
    endcase
  /* decoder.vhd:1979:11  */
  always @*
    case (n4128_o)
      2'b10: n4137_o = 1'b1;
      2'b01: n4137_o = 1'b0;
      default: n4137_o = 1'b0;
    endcase
  /* decoder.vhd:1979:11  */
  always @*
    case (n4128_o)
      2'b10: n4140_o = 4'b0010;
      2'b01: n4140_o = 4'b1100;
      default: n4140_o = 4'b1100;
    endcase
  /* decoder.vhd:1978:9  */
  assign n4142_o = clk_second_cycle_i ? n4131_o : 1'b0;
  /* decoder.vhd:1978:9  */
  assign n4144_o = clk_second_cycle_i ? n4134_o : 1'b0;
  /* decoder.vhd:1978:9  */
  assign n4146_o = clk_second_cycle_i ? n4137_o : 1'b0;
  /* decoder.vhd:1978:9  */
  assign n4148_o = clk_second_cycle_i ? n4140_o : 4'b1100;
  /* decoder.vhd:1975:7  */
  assign n4150_o = opc_mnemonic_s == 6'b111001;
  assign n4151_o = {n4150_o, n4120_o, n4070_o, n4014_o, n4004_o, n3989_o, n3982_o, n3972_o, n3957_o, n3928_o, n3900_o, n3828_o, n3792_o, n3782_o, n3670_o, n3640_o, n3590_o, n3588_o, n3522_o, n3491_o, n3426_o, n3358_o, n3333_o, n3323_o, n3289_o, n3254_o, n3241_o, n3228_o, n3189_o, n3181_o, n3145_o, n3114_o, n3078_o, n3052_o, n3026_o, n3000_o, n2973_o, n2942_o, n2908_o, n2877_o, n2846_o, n2785_o, n2774_o, n2764_o, n2744_o, n2737_o, n2721_o, n2657_o, n2642_o, n2627_o, n2591_o, n2545_o, n2524_o, n2514_o, n2501_o, n2485_o, n2478_o, n2465_o, n2347_o, n2235_o, n2205_o, n2155_o, n2103_o};
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4153_o = n4142_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4153_o = n4103_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4153_o = n4049_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4153_o = n4009_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4153_o = n3943_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4153_o = n3914_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4153_o = n3662_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4153_o = n3623_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4153_o = n3577_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4153_o = n3514_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4153_o = n3479_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4153_o = n3350_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4153_o = n3233_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4153_o = n3217_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4153_o = n3187_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4153_o = n2829_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4153_o = n2780_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4153_o = n2769_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4153_o = n2758_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4153_o = n2613_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4153_o = n2567_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4153_o = n2506_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4153_o = n2470_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4153_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4153_o = n2227_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4153_o = n2188_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4153_o = n2139_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4153_o = n2076_o;
      default: n4153_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4156_o = n3758_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4156_o = n2831_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4156_o = n2701_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4156_o = n2615_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4156_o = n2569_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4156_o = n2323_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4156_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4156_o = 1'b0;
      default: n4156_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4159_o = n4144_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4159_o = n4106_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4159_o = n4052_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4159_o = n3760_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4159_o = n3664_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4159_o = n3626_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4159_o = n3220_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4159_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4159_o = n2325_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4159_o = n2229_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4159_o = n2191_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4159_o = n2141_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4159_o = n2079_o;
      default: n4159_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4162_o = n4146_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4162_o = n4109_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4162_o = n4055_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4162_o = n4012_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4162_o = n3946_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4162_o = n3917_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4162_o = n3820_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4162_o = n3787_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4162_o = n3762_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4162_o = n3666_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4162_o = n3629_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4162_o = n3578_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4162_o = n3516_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4162_o = n3418_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4162_o = n3352_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4162_o = n3328_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4162_o = n3279_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4162_o = n3246_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4162_o = n3171_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4162_o = n2992_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4162_o = n2869_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4162_o = n2834_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4162_o = n2703_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4162_o = n2618_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4162_o = n2572_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4162_o = n2509_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4162_o = n2473_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4162_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4162_o = n2327_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4162_o = n2231_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4162_o = n2194_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4162_o = n2143_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4162_o = n2082_o;
      default: n4162_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4165_o = n3822_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4165_o = n3790_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4165_o = n3764_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4165_o = n3579_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4165_o = n2329_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4165_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4165_o = 1'b0;
      default: n4165_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4168_o = n2436_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4168_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4168_o = 1'b0;
      default: n4168_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4171_o = n2733_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4171_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4171_o = 1'b0;
      default: n4171_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4174_o = n2735_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4174_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4174_o = 1'b0;
      default: n4174_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4177_o = n3331_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4177_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4177_o = 1'b0;
      default: n4177_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4179_o = n4110_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4179_o = n4056_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4179_o = n3881_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4179_o = n3630_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4179_o = n3304_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4179_o = n3280_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4179_o = n3221_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4179_o = n2835_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4179_o = n2437_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4179_o = n2195_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4179_o = n2030_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4179_o = n2083_o;
      default: n4179_o = n2030_o;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4181_o = n4113_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4181_o = n4059_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4181_o = n3882_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4181_o = n3633_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4181_o = n3581_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4181_o = n3313_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4181_o = n3282_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4181_o = n3224_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4181_o = n2837_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4181_o = n2705_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4181_o = n2620_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4181_o = n2198_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4181_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4181_o = n2086_o;
      default: n4181_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4184_o = n3824_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4184_o = n3766_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4184_o = n2331_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4184_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4184_o = 1'b0;
      default: n4184_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4187_o = n3768_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4187_o = n2760_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4187_o = n2333_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4187_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4187_o = 1'b0;
      default: n4187_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4190_o = n3826_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4190_o = n3770_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4190_o = n2335_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4190_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4190_o = 1'b0;
      default: n4190_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4193_o = n3481_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4193_o = n3420_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4193_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4193_o = 1'b0;
      default: n4193_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4196_o = n3772_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4196_o = n3483_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4196_o = n2762_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4196_o = n2337_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4196_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4196_o = 1'b0;
      default: n4196_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4199_o = n3485_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4199_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4199_o = 1'b0;
      default: n4199_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4202_o = n3884_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4202_o = n3173_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4202_o = n3137_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4202_o = n3106_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4202_o = n3072_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4202_o = n3046_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4202_o = n3020_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4202_o = n2994_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4202_o = n2965_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4202_o = n2934_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4202_o = n2900_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4202_o = n2871_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4202_o = n2707_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4202_o = n2439_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4202_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4202_o = 1'b0;
      default: n4202_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4205_o = n2441_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4205_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4205_o = 1'b0;
      default: n4205_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4208_o = n3886_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4208_o = n2967_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4208_o = n2443_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4208_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4208_o = 1'b0;
      default: n4208_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4211_o = n2445_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4211_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4211_o = 1'b0;
      default: n4211_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4214_o = n3236_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4214_o = n2447_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4214_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4214_o = 1'b0;
      default: n4214_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4217_o = n3888_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4217_o = n3239_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4217_o = n2449_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4217_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4217_o = 1'b0;
      default: n4217_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4220_o = n3890_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4220_o = n3249_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4220_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4220_o = 1'b0;
      default: n4220_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4223_o = n3252_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4223_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4223_o = 1'b0;
      default: n4223_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4227_o = n4148_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4227_o = n4116_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4227_o = n4061_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4227_o = 4'b0111;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4227_o = n3949_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4227_o = n3920_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4227_o = n3774_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4227_o = n3668_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4227_o = n3636_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4227_o = n2840_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4227_o = n2709_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4227_o = n2623_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4227_o = n2574_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4227_o = n2512_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4227_o = n2476_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4227_o = 4'b1100;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4227_o = n2339_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4227_o = n2233_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4227_o = n2201_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4227_o = n2145_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4227_o = n2089_o;
      default: n4227_o = 4'b1100;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4230_o = n3951_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4230_o = n3922_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4230_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4230_o = n2147_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4230_o = n2091_o;
      default: n4230_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4233_o = n2578_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4233_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4233_o = 1'b0;
      default: n4233_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4236_o = n4063_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4236_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4236_o = 1'b0;
      default: n4236_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4239_o = n2581_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4239_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4239_o = 1'b0;
      default: n4239_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4242_o = n2584_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4242_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4242_o = 1'b0;
      default: n4242_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4246_o = 1'b1;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4246_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4246_o = 1'b0;
      default: n4246_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4251_o = 1'b1;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4251_o = 1'b1;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4251_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4251_o = 1'b0;
      default: n4251_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4255_o = n3527_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4255_o = 1'b1;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4255_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4255_o = 1'b0;
      default: n4255_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4258_o = n3797_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4258_o = n3530_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4258_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4258_o = 1'b0;
      default: n4258_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4261_o = n3175_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4261_o = n3139_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4261_o = n3108_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4261_o = n3074_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4261_o = n3048_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4261_o = n3022_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4261_o = n2936_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4261_o = n2902_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4261_o = n2873_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4261_o = n2711_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4261_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4261_o = 1'b0;
      default: n4261_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4271_o = 4'b0001;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4271_o = 4'b1000;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4271_o = n3083_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4271_o = 4'b1010;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4271_o = 4'b1001;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4271_o = 4'b0101;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4271_o = n2938_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4271_o = 4'b0010;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4271_o = n2713_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4271_o = 4'b0000;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4271_o = 4'b0000;
      default: n4271_o = 4'b0000;
    endcase
  assign n4273_o = opc_opcode_q[5];
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4274_o = n3157_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4274_o = n3092_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4274_o = n2886_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4274_o = n2715_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4274_o = n4273_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4274_o = n4273_o;
      default: n4274_o = n4273_o;
    endcase
  assign n4275_o = opc_opcode_q[7:6];
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4277_o = n4118_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4277_o = n4065_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4277_o = n3892_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4277_o = n3638_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4277_o = n3315_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4277_o = n3284_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4277_o = n3226_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4277_o = n2842_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4277_o = n2451_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4277_o = n2203_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4277_o = 2'b01;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4277_o = n2093_o;
      default: n4277_o = 2'b01;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4280_o = n3776_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4280_o = n2341_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4280_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4280_o = 1'b0;
      default: n4280_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4283_o = n3778_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4283_o = n2343_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4283_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4283_o = 1'b0;
      default: n4283_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4286_o = n3518_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4286_o = n2996_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4286_o = 2'b00;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4286_o = 2'b00;
      default: n4286_o = 2'b00;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4289_o = n3977_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4289_o = n3953_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4289_o = n3924_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4289_o = n2586_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4289_o = n2539_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4289_o = n2519_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4289_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4289_o = n2149_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4289_o = n2095_o;
      default: n4289_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4292_o = n2453_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4292_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4292_o = 1'b0;
      default: n4292_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4295_o = n3894_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4295_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4295_o = 1'b0;
      default: n4295_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4298_o = n3955_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4298_o = n3926_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4298_o = n2589_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4298_o = n2522_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4298_o = n2483_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4298_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4298_o = n2151_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4298_o = n2098_o;
      default: n4298_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4301_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4301_o = n2153_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4301_o = n2101_o;
      default: n4301_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4304_o = n2541_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4304_o = n2497_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4304_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4304_o = 1'b0;
      default: n4304_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4307_o = n3980_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4307_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4307_o = 1'b0;
      default: n4307_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4310_o = n3354_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4310_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4310_o = 1'b0;
      default: n4310_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4313_o = n3356_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4313_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4313_o = 1'b0;
      default: n4313_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4316_o = n4000_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4316_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4316_o = 1'b0;
      default: n4316_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4319_o = n4002_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4319_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4319_o = 1'b0;
      default: n4319_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4322_o = n3987_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4322_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4322_o = 1'b0;
      default: n4322_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4347_o = 1'b1;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4347_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4347_o = 1'b1;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4347_o = 1'b0;
      default: n4347_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4350_o = n3520_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4350_o = n3179_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4350_o = n3141_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4350_o = n3112_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4350_o = n3076_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4350_o = n3050_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4350_o = n3024_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4350_o = n2998_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4350_o = n2969_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4350_o = n2940_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4350_o = n2906_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4350_o = n2875_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4350_o = n2717_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4350_o = n2455_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4350_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4350_o = 1'b0;
      default: n4350_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4353_o = n2457_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4353_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4353_o = 1'b0;
      default: n4353_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4356_o = n3896_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4356_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4356_o = 1'b0;
      default: n4356_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4359_o = n2499_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4359_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4359_o = 1'b0;
      default: n4359_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4362_o = n2543_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4362_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4362_o = 1'b0;
      default: n4362_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4365_o = n3968_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4365_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4365_o = 1'b0;
      default: n4365_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4368_o = n3970_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4368_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4368_o = 1'b0;
      default: n4368_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4371_o = n2742_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4371_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4371_o = 1'b0;
      default: n4371_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4373_o = n3487_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4373_o = n3422_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4373_o = n2970_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4373_o = n2458_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4373_o = n2034_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4373_o = n2034_o;
      default: n4373_o = n2034_o;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4374_o = n3488_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4374_o = n3423_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4374_o = n2971_o;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4374_o = n2459_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4374_o = n2038_o;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4374_o = n2038_o;
      default: n4374_o = n2038_o;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4376_o = n3780_o;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4376_o = n3583_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4376_o = n2783_o;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4376_o = n2772_o;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4376_o = n2345_o;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4376_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4376_o = 1'b0;
      default: n4376_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4379_o = n4068_o;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4379_o = n3321_o;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4379_o = n3287_o;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4379_o = n2844_o;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4379_o = n2719_o;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4379_o = n2625_o;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4379_o = n2461_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4379_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4379_o = 1'b0;
      default: n4379_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4382_o = n3489_o;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4382_o = n3424_o;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4382_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4382_o = 1'b0;
      default: n4382_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4385_o = n3586_o;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4385_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4385_o = 1'b0;
      default: n4385_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4388_o = n3143_o;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4388_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4388_o = 1'b0;
      default: n4388_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4391_o = n2653_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4391_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4391_o = 1'b0;
      default: n4391_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4394_o = n2655_o;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4394_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4394_o = 1'b0;
      default: n4394_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4397_o = n2638_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4397_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4397_o = 1'b0;
      default: n4397_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4400_o = n2640_o;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4400_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4400_o = 1'b0;
      default: n4400_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4403_o = n3898_o;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4403_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4403_o = 1'b0;
      default: n4403_o = 1'b0;
    endcase
  /* decoder.vhd:635:5  */
  always @*
    case (n4151_o)
      63'b100000000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b010000000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b001000000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000100000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000010000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000001000000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000100000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000010000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000001000000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000100000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000010000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000001000000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000100000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000010000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000001000000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000100000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000010000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000001000000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000100000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000010000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000001000000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000100000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000010000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000001000000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000100000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000010000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000001000000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000100000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000010000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000001000000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000100000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000010000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000001000000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000100000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000010000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000001000000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000100000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000010000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000001000000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000100000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000010000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000001000000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000100000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000010000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000001000000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000100000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000010000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000001000000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000100000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000010000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000001000000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000100000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000010000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000001000000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000100000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000010000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000001000000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000100000: n4406_o = n2463_o;
      63'b000000000000000000000000000000000000000000000000000000000010000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000001000: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000100: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000010: n4406_o = 1'b0;
      63'b000000000000000000000000000000000000000000000000000000000000001: n4406_o = 1'b0;
      default: n4406_o = 1'b0;
    endcase
  /* decoder.vhd:2020:14  */
  assign n4410_o = ~res_i;
  /* decoder.vhd:2035:7  */
  assign n4413_o = bus_clear_f1_i ? 1'b0 : f1_q;
  /* decoder.vhd:2033:7  */
  assign n4415_o = bus_set_f1_i ? 1'b1 : n4413_o;
  /* decoder.vhd:2044:28  */
  assign n4417_o = clk_mstate_i == 3'b100;
  /* decoder.vhd:2044:9  */
  assign n4419_o = n4417_o ? 1'b0 : branch_taken_q;
  /* decoder.vhd:2042:9  */
  assign n4421_o = branch_taken_s ? 1'b1 : n4419_o;
  /* decoder.vhd:2053:27  */
  assign n4422_o = ~f1_q;
  /* decoder.vhd:2052:9  */
  assign n4423_o = cpl_f1_s ? n4422_o : n4415_o;
  /* decoder.vhd:2050:9  */
  assign n4425_o = clear_f1_s ? 1'b0 : n4423_o;
  /* decoder.vhd:2059:9  */
  assign n4427_o = set_mb_s ? 1'b1 : mb_q;
  /* decoder.vhd:2057:9  */
  assign n4429_o = clear_mb_s ? 1'b0 : n4427_o;
  /* decoder.vhd:2039:7  */
  assign n4433_o = en_clk_i ? n4425_o : n4415_o;
  /* decoder.vhd:2039:7  */
  assign n4435_o = en_clk_i & ent0_clk_s;
  /* decoder.vhd:2115:27  */
  assign n4449_o = read_dec_s ? data_s : 8'b11111111;
  /* decoder.vhd:2117:48  */
  assign n4451_o = en_clk_i & dm_write_dmem_s;
  /* decoder.vhd:2118:48  */
  assign n4452_o = pm_inc_pc_s | add_inc_pc_s;
  /* decoder.vhd:2119:48  */
  assign n4453_o = pm_write_pmem_addr_s | add_write_pmem_addr_s;
  /* decoder.vhd:2121:48  */
  assign n4454_o = bus_read_bus_s | add_read_bus_s;
  /* decoder.vhd:305:5  */
  assign n4455_o = en_clk_i ? n1869_o : opc_opcode_q;
  /* decoder.vhd:305:5  */
  always @(posedge clk_i or posedge n1863_o)
    if (n1863_o)
      n4456_q <= 8'b00000000;
    else
      n4456_q <= n4455_o;
  /* decoder.vhd:2031:5  */
  assign n4457_o = en_clk_i ? n4421_o : branch_taken_q;
  /* decoder.vhd:2031:5  */
  always @(posedge clk_i or posedge n4410_o)
    if (n4410_o)
      n4458_q <= 1'b0;
    else
      n4458_q <= n4457_o;
  /* decoder.vhd:2031:5  */
  always @(posedge clk_i or posedge n4410_o)
    if (n4410_o)
      n4459_q <= 1'b0;
    else
      n4459_q <= n4433_o;
  /* decoder.vhd:2031:5  */
  assign n4460_o = en_clk_i ? n4429_o : mb_q;
  /* decoder.vhd:2031:5  */
  always @(posedge clk_i or posedge n4410_o)
    if (n4410_o)
      n4461_q <= 1'b0;
    else
      n4461_q <= n4460_o;
  /* decoder.vhd:2031:5  */
  assign n4462_o = n4435_o ? 1'b1 : t0_dir_q;
  /* decoder.vhd:2031:5  */
  always @(posedge clk_i or posedge n4410_o)
    if (n4410_o)
      n4463_q <= 1'b0;
    else
      n4463_q <= n4462_o;
  /* decoder.vhd:305:5  */
  assign n4464_o = en_clk_i ? n1870_o : mnemonic_q;
  /* decoder.vhd:305:5  */
  always @(posedge clk_i or posedge n1863_o)
    if (n1863_o)
      n4465_q <= 6'b101001;
    else
      n4465_q <= n4464_o;
  /* decoder.vhd:301:5  */
  assign n4466_o = {n4275_o, n4274_o};
endmodule

module t48_db_bus
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  ea_i,
   input  [7:0] data_i,
   input  write_bus_i,
   input  read_bus_i,
   input  output_pcl_i,
   input  bidir_bus_i,
   input  [7:0] pcl_i,
   input  [7:0] db_i,
   output [7:0] data_o,
   output [7:0] db_o,
   output db_dir_o);
  wire [7:0] bus_q;
  wire db_dir_q;
  wire db_dir_qq;
  wire n998_o;
  wire n1001_o;
  wire n1002_o;
  wire n1004_o;
  wire n1007_o;
  wire n1008_o;
  wire [7:0] n1021_o;
  wire n1029_o;
  wire n1030_o;
  wire n1032_o;
  wire [7:0] n1033_o;
  wire [7:0] n1034_o;
  reg [7:0] n1035_q;
  wire n1036_o;
  reg n1037_q;
  wire n1038_o;
  reg n1039_q;
  assign data_o = n1033_o;
  assign db_o = n1021_o;
  assign db_dir_o = n1030_o;
  /* db_bus.vhd:85:10  */
  assign bus_q = n1035_q; // (signal)
  /* db_bus.vhd:88:10  */
  assign db_dir_q = n1037_q; // (signal)
  /* db_bus.vhd:89:10  */
  assign db_dir_qq = n1039_q; // (signal)
  /* db_bus.vhd:101:14  */
  assign n998_o = ~res_i;
  /* db_bus.vhd:108:9  */
  assign n1001_o = write_bus_i ? 1'b1 : db_dir_q;
  /* db_bus.vhd:120:26  */
  assign n1002_o = ea_i | bidir_bus_i;
  /* db_bus.vhd:120:9  */
  assign n1004_o = n1002_o ? 1'b0 : db_dir_q;
  /* db_bus.vhd:115:9  */
  assign n1007_o = write_bus_i ? 1'b1 : n1004_o;
  /* db_bus.vhd:107:7  */
  assign n1008_o = en_clk_i & write_bus_i;
  /* db_bus.vhd:138:15  */
  assign n1021_o = output_pcl_i ? pcl_i : bus_q;
  /* t48_pack-p.vhd:66:5  */
  assign n1029_o = output_pcl_i ? 1'b1 : 1'b0;
  /* db_bus.vhd:140:25  */
  assign n1030_o = db_dir_qq | n1029_o;
  /* db_bus.vhd:143:20  */
  assign n1032_o = ~read_bus_i;
  /* db_bus.vhd:143:15  */
  assign n1033_o = n1032_o ? 8'b11111111 : db_i;
  /* db_bus.vhd:106:5  */
  assign n1034_o = n1008_o ? data_i : bus_q;
  /* db_bus.vhd:106:5  */
  always @(posedge clk_i or posedge n998_o)
    if (n998_o)
      n1035_q <= 8'b00000000;
    else
      n1035_q <= n1034_o;
  /* db_bus.vhd:106:5  */
  assign n1036_o = en_clk_i ? n1007_o : db_dir_q;
  /* db_bus.vhd:106:5  */
  always @(posedge clk_i or posedge n998_o)
    if (n998_o)
      n1037_q <= 1'b0;
    else
      n1037_q <= n1036_o;
  /* db_bus.vhd:106:5  */
  assign n1038_o = en_clk_i ? n1001_o : db_dir_qq;
  /* db_bus.vhd:106:5  */
  always @(posedge clk_i or posedge n998_o)
    if (n998_o)
      n1039_q <= 1'b0;
    else
      n1039_q <= n1038_o;
endmodule

module t48_cond_branch
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  compute_take_i,
   input  [3:0] branch_cond_i,
   input  [7:0] accu_i,
   input  t0_i,
   input  t1_i,
   input  int_n_i,
   input  f0_i,
   input  f1_i,
   input  tf_i,
   input  carry_i,
   input  ibf_i,
   input  obf_i,
   input  [2:0] comp_value_i,
   output take_branch_o);
  wire take_branch_s;
  wire take_branch_q;
  wire n910_o;
  wire n912_o;
  wire n913_o;
  wire n915_o;
  wire n916_o;
  wire n917_o;
  wire n918_o;
  wire n919_o;
  wire n920_o;
  wire n921_o;
  wire n922_o;
  wire n923_o;
  wire n924_o;
  wire n925_o;
  wire n926_o;
  wire n927_o;
  wire n928_o;
  wire n929_o;
  wire n930_o;
  wire n931_o;
  wire n932_o;
  wire n934_o;
  wire n935_o;
  wire n936_o;
  wire n938_o;
  wire n940_o;
  wire n942_o;
  wire n943_o;
  wire n945_o;
  wire n946_o;
  wire n947_o;
  wire n949_o;
  wire n950_o;
  wire n951_o;
  wire n953_o;
  wire n955_o;
  wire n956_o;
  wire n958_o;
  wire n960_o;
  wire [10:0] n961_o;
  reg n963_o;
  wire n970_o;
  wire n973_o;
  wire n978_o;
  reg n979_q;
  wire n980_o;
  wire n981_o;
  wire n982_o;
  wire n983_o;
  wire n984_o;
  wire n985_o;
  wire n986_o;
  wire n987_o;
  wire [1:0] n988_o;
  reg n989_o;
  wire [1:0] n990_o;
  reg n991_o;
  wire n992_o;
  wire n993_o;
  assign take_branch_o = take_branch_q;
  /* cond_branch.vhd:90:10  */
  assign take_branch_s = n963_o; // (signal)
  /* cond_branch.vhd:91:10  */
  assign take_branch_q = n979_q; // (signal)
  /* cond_branch.vhd:119:9  */
  assign n910_o = n993_o ? 1'b1 : 1'b0;
  /* cond_branch.vhd:118:7  */
  assign n912_o = branch_cond_i == 4'b0000;
  /* cond_branch.vhd:126:33  */
  assign n913_o = accu_i[7];
  /* cond_branch.vhd:126:24  */
  assign n915_o = 1'b0 | n913_o;
  /* cond_branch.vhd:126:33  */
  assign n916_o = accu_i[6];
  /* cond_branch.vhd:126:24  */
  assign n917_o = n915_o | n916_o;
  /* cond_branch.vhd:126:33  */
  assign n918_o = accu_i[5];
  /* cond_branch.vhd:126:24  */
  assign n919_o = n917_o | n918_o;
  /* cond_branch.vhd:126:33  */
  assign n920_o = accu_i[4];
  /* cond_branch.vhd:126:24  */
  assign n921_o = n919_o | n920_o;
  /* cond_branch.vhd:126:33  */
  assign n922_o = accu_i[3];
  /* cond_branch.vhd:126:24  */
  assign n923_o = n921_o | n922_o;
  /* cond_branch.vhd:126:33  */
  assign n924_o = accu_i[2];
  /* cond_branch.vhd:126:24  */
  assign n925_o = n923_o | n924_o;
  /* cond_branch.vhd:126:33  */
  assign n926_o = accu_i[1];
  /* cond_branch.vhd:126:24  */
  assign n927_o = n925_o | n926_o;
  /* cond_branch.vhd:126:33  */
  assign n928_o = accu_i[0];
  /* cond_branch.vhd:126:24  */
  assign n929_o = n927_o | n928_o;
  /* cond_branch.vhd:128:49  */
  assign n930_o = comp_value_i[0];
  /* cond_branch.vhd:128:33  */
  assign n931_o = ~n930_o;
  /* cond_branch.vhd:128:31  */
  assign n932_o = n929_o == n931_o;
  /* cond_branch.vhd:124:7  */
  assign n934_o = branch_cond_i == 4'b0001;
  /* cond_branch.vhd:132:48  */
  assign n935_o = comp_value_i[0];
  /* cond_branch.vhd:132:34  */
  assign n936_o = carry_i == n935_o;
  /* cond_branch.vhd:131:7  */
  assign n938_o = branch_cond_i == 4'b0010;
  /* cond_branch.vhd:135:7  */
  assign n940_o = branch_cond_i == 4'b0011;
  /* cond_branch.vhd:139:7  */
  assign n942_o = branch_cond_i == 4'b0100;
  /* cond_branch.vhd:144:34  */
  assign n943_o = ~int_n_i;
  /* cond_branch.vhd:143:7  */
  assign n945_o = branch_cond_i == 4'b0101;
  /* cond_branch.vhd:148:45  */
  assign n946_o = comp_value_i[0];
  /* cond_branch.vhd:148:31  */
  assign n947_o = t0_i == n946_o;
  /* cond_branch.vhd:147:7  */
  assign n949_o = branch_cond_i == 4'b0110;
  /* cond_branch.vhd:152:45  */
  assign n950_o = comp_value_i[0];
  /* cond_branch.vhd:152:31  */
  assign n951_o = t1_i == n950_o;
  /* cond_branch.vhd:151:7  */
  assign n953_o = branch_cond_i == 4'b0111;
  /* cond_branch.vhd:155:7  */
  assign n955_o = branch_cond_i == 4'b1000;
  /* cond_branch.vhd:160:32  */
  assign n956_o = ~ibf_i;
  /* cond_branch.vhd:159:7  */
  assign n958_o = branch_cond_i == 4'b1001;
  /* cond_branch.vhd:163:7  */
  assign n960_o = branch_cond_i == 4'b1010;
  /* clock_ctrl.vhd:206:5  */
  assign n961_o = {n960_o, n958_o, n955_o, n953_o, n949_o, n945_o, n942_o, n940_o, n938_o, n934_o, n912_o};
  /* cond_branch.vhd:116:5  */
  always @*
    case (n961_o)
      11'b10000000000: n963_o = obf_i;
      11'b01000000000: n963_o = n956_o;
      11'b00100000000: n963_o = tf_i;
      11'b00010000000: n963_o = n951_o;
      11'b00001000000: n963_o = n947_o;
      11'b00000100000: n963_o = n943_o;
      11'b00000010000: n963_o = f1_i;
      11'b00000001000: n963_o = f0_i;
      11'b00000000100: n963_o = n936_o;
      11'b00000000010: n963_o = n932_o;
      11'b00000000001: n963_o = n910_o;
      default: n963_o = 1'b0;
    endcase
  /* cond_branch.vhd:188:14  */
  assign n970_o = ~res_i;
  /* cond_branch.vhd:192:7  */
  assign n973_o = en_clk_i & compute_take_i;
  /* cond_branch.vhd:191:5  */
  assign n978_o = n973_o ? take_branch_s : take_branch_q;
  /* cond_branch.vhd:191:5  */
  always @(posedge clk_i or posedge n970_o)
    if (n970_o)
      n979_q <= 1'b0;
    else
      n979_q <= n978_o;
  /* cond_branch.vhd:64:5  */
  assign n980_o = accu_i[0];
  assign n981_o = accu_i[1];
  /* cond_branch.vhd:191:5  */
  assign n982_o = accu_i[2];
  /* cond_branch.vhd:186:3  */
  assign n983_o = accu_i[3];
  assign n984_o = accu_i[4];
  assign n985_o = accu_i[5];
  /* cond_branch.vhd:116:5  */
  assign n986_o = accu_i[6];
  assign n987_o = accu_i[7];
  /* cond_branch.vhd:119:18  */
  assign n988_o = comp_value_i[1:0];
  /* cond_branch.vhd:119:18  */
  always @*
    case (n988_o)
      2'b00: n989_o = n980_o;
      2'b01: n989_o = n981_o;
      2'b10: n989_o = n982_o;
      2'b11: n989_o = n983_o;
    endcase
  /* cond_branch.vhd:119:18  */
  assign n990_o = comp_value_i[1:0];
  /* cond_branch.vhd:119:18  */
  always @*
    case (n990_o)
      2'b00: n991_o = n984_o;
      2'b01: n991_o = n985_o;
      2'b10: n991_o = n986_o;
      2'b11: n991_o = n987_o;
    endcase
  /* cond_branch.vhd:119:18  */
  assign n992_o = comp_value_i[2];
  /* cond_branch.vhd:119:18  */
  assign n993_o = n992_o ? n991_o : n989_o;
endmodule

module t48_clock_ctrl_1
  (input  clk_i,
   input  xtal_i,
   input  xtal_en_i,
   input  res_i,
   input  en_clk_i,
   input  multi_cycle_i,
   input  assert_psen_i,
   input  assert_prog_i,
   input  assert_rd_i,
   input  assert_wr_i,
   output xtal3_o,
   output t0_o,
   output [2:0] mstate_o,
   output second_cycle_o,
   output ale_o,
   output psen_o,
   output prog_o,
   output rd_o,
   output wr_o);
  wire [1:0] xtal_q;
  wire xtal2_s;
  wire xtal3_s;
  wire x2_s;
  wire x3_s;
  wire t0_q;
  wire [2:0] mstate_q;
  wire ale_q;
  wire psen_q;
  wire prog_q;
  wire rd_q;
  wire wr_q;
  wire second_cycle_q;
  wire multi_cycle_q;
  wire n686_o;
  wire n689_o;
  wire [1:0] n691_o;
  wire [1:0] n693_o;
  wire n696_o;
  wire n714_o;
  wire n715_o;
  wire n716_o;
  wire n720_o;
  wire n721_o;
  wire n722_o;
  wire n739_o;
  wire n747_o;
  wire n749_o;
  wire n751_o;
  wire n752_o;
  wire n754_o;
  wire n756_o;
  wire n757_o;
  wire n758_o;
  wire n760_o;
  wire n762_o;
  wire n764_o;
  wire n766_o;
  wire n768_o;
  wire n770_o;
  wire n772_o;
  wire n774_o;
  wire n776_o;
  wire n778_o;
  wire n779_o;
  wire n780_o;
  wire n781_o;
  wire n782_o;
  wire n783_o;
  wire n785_o;
  wire n787_o;
  wire n789_o;
  wire [4:0] n790_o;
  reg n792_o;
  reg n794_o;
  reg n796_o;
  reg n798_o;
  reg n800_o;
  wire n818_o;
  wire n821_o;
  wire n823_o;
  wire n825_o;
  wire n827_o;
  wire n829_o;
  wire [4:0] n830_o;
  reg [2:0] n837_o;
  wire n846_o;
  wire n849_o;
  wire n851_o;
  wire n852_o;
  wire n854_o;
  wire n855_o;
  wire n857_o;
  wire n858_o;
  wire n859_o;
  wire n861_o;
  wire n863_o;
  wire [1:0] n887_o;
  reg [1:0] n888_q;
  wire n889_o;
  reg n890_q;
  wire [2:0] n891_o;
  reg [2:0] n892_q;
  reg n893_q;
  reg n894_q;
  reg n895_q;
  reg n896_q;
  reg n897_q;
  wire n898_o;
  reg n899_q;
  wire n900_o;
  reg n901_q;
  assign xtal3_o = xtal3_s;
  assign t0_o = t0_q;
  assign mstate_o = mstate_q;
  assign second_cycle_o = second_cycle_q;
  assign ale_o = ale_q;
  assign psen_o = psen_q;
  assign prog_o = prog_q;
  assign rd_o = rd_q;
  assign wr_o = wr_q;
  /* clock_ctrl.vhd:90:10  */
  assign xtal_q = n888_q; // (signal)
  /* clock_ctrl.vhd:92:10  */
  assign xtal2_s = n739_o; // (signal)
  /* clock_ctrl.vhd:93:10  */
  assign xtal3_s = n747_o; // (signal)
  /* clock_ctrl.vhd:95:10  */
  assign x2_s = n716_o; // (signal)
  /* clock_ctrl.vhd:96:10  */
  assign x3_s = n722_o; // (signal)
  /* clock_ctrl.vhd:98:10  */
  assign t0_q = n890_q; // (signal)
  /* clock_ctrl.vhd:102:10  */
  assign mstate_q = n892_q; // (signal)
  /* clock_ctrl.vhd:104:10  */
  assign ale_q = n893_q; // (signal)
  /* clock_ctrl.vhd:105:10  */
  assign psen_q = n894_q; // (signal)
  /* clock_ctrl.vhd:106:10  */
  assign prog_q = n895_q; // (signal)
  /* clock_ctrl.vhd:107:10  */
  assign rd_q = n896_q; // (signal)
  /* clock_ctrl.vhd:108:10  */
  assign wr_q = n897_q; // (signal)
  /* clock_ctrl.vhd:112:10  */
  assign second_cycle_q = n899_q; // (signal)
  /* clock_ctrl.vhd:113:10  */
  assign multi_cycle_q = n901_q; // (signal)
  /* clock_ctrl.vhd:137:16  */
  assign n686_o = ~res_i;
  /* clock_ctrl.vhd:143:21  */
  assign n689_o = $unsigned(xtal_q) < $unsigned(2'b10);
  /* clock_ctrl.vhd:144:30  */
  assign n691_o = xtal_q + 2'b01;
  /* clock_ctrl.vhd:143:11  */
  assign n693_o = n689_o ? n691_o : 2'b00;
  /* clock_ctrl.vhd:149:11  */
  assign n696_o = xtal3_s ? 1'b1 : 1'b0;
  /* clock_ctrl.vhd:164:25  */
  assign n714_o = xtal_q == 2'b01;
  /* clock_ctrl.vhd:164:29  */
  assign n715_o = xtal_en_i & n714_o;
  /* clock_ctrl.vhd:164:13  */
  assign n716_o = n715_o ? 1'b1 : 1'b0;
  /* clock_ctrl.vhd:167:25  */
  assign n720_o = xtal_q == 2'b10;
  /* clock_ctrl.vhd:167:29  */
  assign n721_o = xtal_en_i & n720_o;
  /* clock_ctrl.vhd:167:13  */
  assign n722_o = n721_o ? 1'b1 : 1'b0;
  /* t48_pack-p.vhd:75:5  */
  assign n739_o = x2_s ? 1'b1 : 1'b0;
  /* t48_pack-p.vhd:75:5  */
  assign n747_o = x3_s ? 1'b1 : 1'b0;
  /* clock_ctrl.vhd:206:14  */
  assign n749_o = ~res_i;
  /* clock_ctrl.vhd:218:26  */
  assign n751_o = ~second_cycle_q;
  /* clock_ctrl.vhd:218:22  */
  assign n752_o = n751_o & xtal2_s;
  /* clock_ctrl.vhd:218:11  */
  assign n754_o = n757_o ? 1'b1 : rd_q;
  /* clock_ctrl.vhd:218:11  */
  assign n756_o = n758_o ? 1'b1 : wr_q;
  /* clock_ctrl.vhd:218:11  */
  assign n757_o = n752_o & assert_rd_i;
  /* clock_ctrl.vhd:218:11  */
  assign n758_o = n752_o & assert_wr_i;
  /* clock_ctrl.vhd:216:9  */
  assign n760_o = mstate_q == 3'b100;
  /* clock_ctrl.vhd:228:11  */
  assign n762_o = xtal3_s ? 1'b0 : psen_q;
  /* clock_ctrl.vhd:227:9  */
  assign n764_o = mstate_q == 3'b000;
  /* clock_ctrl.vhd:233:11  */
  assign n766_o = xtal3_s ? 1'b0 : prog_q;
  /* clock_ctrl.vhd:233:11  */
  assign n768_o = xtal3_s ? 1'b0 : rd_q;
  /* clock_ctrl.vhd:233:11  */
  assign n770_o = xtal3_s ? 1'b0 : wr_q;
  /* clock_ctrl.vhd:232:9  */
  assign n772_o = mstate_q == 3'b001;
  /* clock_ctrl.vhd:243:11  */
  assign n774_o = xtal3_s ? 1'b1 : ale_q;
  /* clock_ctrl.vhd:241:9  */
  assign n776_o = mstate_q == 3'b010;
  /* clock_ctrl.vhd:248:11  */
  assign n778_o = n779_o ? 1'b1 : psen_q;
  /* clock_ctrl.vhd:248:11  */
  assign n779_o = xtal3_s & assert_psen_i;
  /* clock_ctrl.vhd:257:22  */
  assign n780_o = multi_cycle_q & xtal3_s;
  /* clock_ctrl.vhd:258:32  */
  assign n781_o = ~second_cycle_q;
  /* clock_ctrl.vhd:258:28  */
  assign n782_o = n781_o & n780_o;
  /* clock_ctrl.vhd:258:51  */
  assign n783_o = assert_prog_i & n782_o;
  /* clock_ctrl.vhd:257:11  */
  assign n785_o = n783_o ? 1'b1 : prog_q;
  /* clock_ctrl.vhd:263:11  */
  assign n787_o = xtal2_s ? 1'b0 : ale_q;
  /* clock_ctrl.vhd:247:9  */
  assign n789_o = mstate_q == 3'b011;
  assign n790_o = {n789_o, n776_o, n772_o, n764_o, n760_o};
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n790_o)
      5'b10000: n792_o = n787_o;
      5'b01000: n792_o = n774_o;
      5'b00100: n792_o = ale_q;
      5'b00010: n792_o = ale_q;
      5'b00001: n792_o = ale_q;
      default: n792_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n790_o)
      5'b10000: n794_o = n778_o;
      5'b01000: n794_o = psen_q;
      5'b00100: n794_o = psen_q;
      5'b00010: n794_o = n762_o;
      5'b00001: n794_o = psen_q;
      default: n794_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n790_o)
      5'b10000: n796_o = n785_o;
      5'b01000: n796_o = prog_q;
      5'b00100: n796_o = n766_o;
      5'b00010: n796_o = prog_q;
      5'b00001: n796_o = prog_q;
      default: n796_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n790_o)
      5'b10000: n798_o = rd_q;
      5'b01000: n798_o = rd_q;
      5'b00100: n798_o = n768_o;
      5'b00010: n798_o = rd_q;
      5'b00001: n798_o = n754_o;
      default: n798_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:215:7  */
  always @*
    case (n790_o)
      5'b10000: n800_o = wr_q;
      5'b01000: n800_o = wr_q;
      5'b00100: n800_o = n770_o;
      5'b00010: n800_o = wr_q;
      5'b00001: n800_o = n756_o;
      default: n800_o = 1'b0;
    endcase
  /* clock_ctrl.vhd:292:14  */
  assign n818_o = ~res_i;
  /* clock_ctrl.vhd:303:11  */
  assign n821_o = mstate_q == 3'b100;
  /* clock_ctrl.vhd:306:11  */
  assign n823_o = mstate_q == 3'b000;
  /* clock_ctrl.vhd:309:11  */
  assign n825_o = mstate_q == 3'b001;
  /* clock_ctrl.vhd:312:11  */
  assign n827_o = mstate_q == 3'b010;
  /* clock_ctrl.vhd:315:11  */
  assign n829_o = mstate_q == 3'b011;
  assign n830_o = {n829_o, n827_o, n825_o, n823_o, n821_o};
  /* clock_ctrl.vhd:302:9  */
  always @*
    case (n830_o)
      5'b10000: n837_o = 3'b100;
      5'b01000: n837_o = 3'b011;
      5'b00100: n837_o = 3'b010;
      5'b00010: n837_o = 3'b001;
      5'b00001: n837_o = 3'b000;
      default: n837_o = 3'b000;
    endcase
  /* clock_ctrl.vhd:349:14  */
  assign n846_o = ~res_i;
  /* clock_ctrl.vhd:356:30  */
  assign n849_o = mstate_q == 3'b001;
  /* clock_ctrl.vhd:357:30  */
  assign n851_o = mstate_q == 3'b100;
  /* clock_ctrl.vhd:360:21  */
  assign n852_o = multi_cycle_i & n849_o;
  /* clock_ctrl.vhd:360:9  */
  assign n854_o = n852_o ? 1'b1 : multi_cycle_q;
  /* clock_ctrl.vhd:365:26  */
  assign n855_o = n851_o & multi_cycle_q;
  /* clock_ctrl.vhd:365:9  */
  assign n857_o = n855_o ? 1'b1 : second_cycle_q;
  /* clock_ctrl.vhd:371:27  */
  assign n858_o = second_cycle_q & multi_cycle_q;
  /* clock_ctrl.vhd:370:21  */
  assign n859_o = n858_o & n851_o;
  /* clock_ctrl.vhd:370:9  */
  assign n861_o = n859_o ? 1'b0 : n857_o;
  /* clock_ctrl.vhd:370:9  */
  assign n863_o = n859_o ? 1'b0 : n854_o;
  /* clock_ctrl.vhd:141:7  */
  assign n887_o = xtal_en_i ? n693_o : xtal_q;
  /* clock_ctrl.vhd:141:7  */
  always @(posedge xtal_i or posedge n686_o)
    if (n686_o)
      n888_q <= 2'b00;
    else
      n888_q <= n887_o;
  /* clock_ctrl.vhd:141:7  */
  assign n889_o = xtal_en_i ? n696_o : t0_q;
  /* clock_ctrl.vhd:141:7  */
  always @(posedge xtal_i or posedge n686_o)
    if (n686_o)
      n890_q <= 1'b0;
    else
      n890_q <= n889_o;
  /* clock_ctrl.vhd:299:5  */
  assign n891_o = en_clk_i ? n837_o : mstate_q;
  /* clock_ctrl.vhd:299:5  */
  always @(posedge clk_i or posedge n818_o)
    if (n818_o)
      n892_q <= 3'b010;
    else
      n892_q <= n891_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n749_o)
    if (n749_o)
      n893_q <= 1'b0;
    else
      n893_q <= n792_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n749_o)
    if (n749_o)
      n894_q <= 1'b0;
    else
      n894_q <= n794_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n749_o)
    if (n749_o)
      n895_q <= 1'b0;
    else
      n895_q <= n796_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n749_o)
    if (n749_o)
      n896_q <= 1'b0;
    else
      n896_q <= n798_o;
  /* clock_ctrl.vhd:213:5  */
  always @(posedge xtal_i or posedge n749_o)
    if (n749_o)
      n897_q <= 1'b0;
    else
      n897_q <= n800_o;
  /* clock_ctrl.vhd:353:5  */
  assign n898_o = en_clk_i ? n861_o : second_cycle_q;
  /* clock_ctrl.vhd:353:5  */
  always @(posedge clk_i or posedge n846_o)
    if (n846_o)
      n899_q <= 1'b0;
    else
      n899_q <= n898_o;
  /* clock_ctrl.vhd:353:5  */
  assign n900_o = en_clk_i ? n863_o : multi_cycle_q;
  /* clock_ctrl.vhd:353:5  */
  always @(posedge clk_i or posedge n846_o)
    if (n846_o)
      n901_q <= 1'b0;
    else
      n901_q <= n900_o;
endmodule

module t48_bus_mux
  (input  [7:0] alu_data_i,
   input  [7:0] bus_data_i,
   input  [7:0] dec_data_i,
   input  [7:0] dm_data_i,
   input  [7:0] pm_data_i,
   input  [7:0] p1_data_i,
   input  [7:0] p2_data_i,
   input  [7:0] psw_data_i,
   input  [7:0] tim_data_i,
   output [7:0] data_o);
  wire [7:0] n668_o;
  wire [7:0] n669_o;
  wire [7:0] n670_o;
  wire [7:0] n671_o;
  wire [7:0] n672_o;
  wire [7:0] n673_o;
  wire [7:0] n674_o;
  wire [7:0] n675_o;
  assign data_o = n675_o;
  /* bus_mux.vhd:89:26  */
  assign n668_o = alu_data_i & bus_data_i;
  /* bus_mux.vhd:90:26  */
  assign n669_o = n668_o & dec_data_i;
  /* bus_mux.vhd:91:26  */
  assign n670_o = n669_o & dm_data_i;
  /* bus_mux.vhd:92:26  */
  assign n671_o = n670_o & pm_data_i;
  /* bus_mux.vhd:93:26  */
  assign n672_o = n671_o & p1_data_i;
  /* bus_mux.vhd:94:26  */
  assign n673_o = n672_o & p2_data_i;
  /* bus_mux.vhd:95:26  */
  assign n674_o = n673_o & psw_data_i;
  /* bus_mux.vhd:96:26  */
  assign n675_o = n674_o & tim_data_i;
endmodule

module t48_alu
  (input  clk_i,
   input  res_i,
   input  en_clk_i,
   input  [7:0] data_i,
   input  write_accu_i,
   input  write_shadow_i,
   input  write_temp_reg_i,
   input  read_alu_i,
   input  carry_i,
   input  [3:0] alu_op_i,
   input  use_carry_i,
   input  da_high_i,
   input  accu_low_i,
   input  p06_temp_reg_i,
   input  p60_temp_reg_i,
   output [7:0] data_o,
   output carry_o,
   output aux_carry_o,
   output da_overflow_o);
  wire [7:0] accumulator_q;
  wire [7:0] accu_shadow_q;
  wire [7:0] temp_req_q;
  wire [7:0] in_a_s;
  wire [7:0] in_b_s;
  wire [7:0] data_s;
  wire [8:0] add_result_s;
  wire n417_o;
  wire [3:0] n419_o;
  wire [3:0] n420_o;
  wire [3:0] n421_o;
  wire [3:0] n422_o;
  wire [3:0] n423_o;
  wire [3:0] n424_o;
  wire [7:0] n425_o;
  wire [7:0] n427_o;
  wire [7:0] n428_o;
  wire [7:0] n430_o;
  wire [7:0] n432_o;
  wire n433_o;
  wire [7:0] n447_o;
  wire n449_o;
  wire [7:0] n450_o;
  wire n452_o;
  wire [7:0] n453_o;
  wire n455_o;
  wire [7:0] n456_o;
  wire n457_o;
  wire n459_o;
  wire [7:0] n460_o;
  wire n462_o;
  wire n464_o;
  wire [6:0] n465_o;
  wire n466_o;
  wire n467_o;
  wire n468_o;
  wire n470_o;
  wire [6:0] n471_o;
  wire n472_o;
  wire n473_o;
  wire n474_o;
  wire n476_o;
  wire [3:0] n477_o;
  wire [3:0] n478_o;
  wire n480_o;
  wire [7:0] n481_o;
  wire n483_o;
  wire [7:0] n484_o;
  wire n486_o;
  wire [3:0] n487_o;
  wire [3:0] n488_o;
  wire [7:0] n489_o;
  wire n491_o;
  wire n493_o;
  wire [12:0] n494_o;
  reg n496_o;
  wire n498_o;
  wire n499_o;
  wire n500_o;
  wire n501_o;
  wire n502_o;
  wire n504_o;
  wire n505_o;
  wire n506_o;
  wire n507_o;
  wire n508_o;
  wire n509_o;
  reg n511_o;
  wire [2:0] n512_o;
  wire [2:0] n513_o;
  wire [2:0] n514_o;
  wire [2:0] n515_o;
  wire [2:0] n516_o;
  wire [2:0] n518_o;
  wire [2:0] n519_o;
  wire [2:0] n520_o;
  wire [2:0] n521_o;
  wire [2:0] n522_o;
  wire [2:0] n523_o;
  wire [2:0] n524_o;
  reg [2:0] n526_o;
  wire [2:0] n527_o;
  wire [2:0] n528_o;
  wire [2:0] n529_o;
  wire [2:0] n530_o;
  wire [2:0] n531_o;
  wire [2:0] n533_o;
  wire [2:0] n534_o;
  wire [2:0] n535_o;
  wire [2:0] n536_o;
  wire [2:0] n537_o;
  wire [2:0] n538_o;
  wire [2:0] n539_o;
  reg [2:0] n541_o;
  wire n542_o;
  wire n543_o;
  wire n544_o;
  wire n545_o;
  wire n546_o;
  wire n548_o;
  wire n549_o;
  wire n550_o;
  wire n551_o;
  wire n552_o;
  wire n553_o;
  reg n555_o;
  wire n567_o;
  wire n570_o;
  localparam [8:0] n571_o = 9'b000000000;
  wire [7:0] n572_o;
  wire [8:0] n574_o;
  wire [8:0] n576_o;
  localparam [8:0] n578_o = 9'b000000000;
  wire [7:0] n579_o;
  wire n581_o;
  wire n583_o;
  wire [1:0] n584_o;
  wire n586_o;
  reg n587_o;
  wire [7:0] n589_o;
  reg [7:0] n590_o;
  wire [8:0] n592_o;
  wire [8:0] n593_o;
  wire [8:0] n594_o;
  wire [8:0] n595_o;
  wire n596_o;
  wire n597_o;
  wire [1:0] n598_o;
  wire n599_o;
  wire n602_o;
  wire n604_o;
  wire n606_o;
  wire n607_o;
  wire n608_o;
  wire n609_o;
  wire n612_o;
  wire n614_o;
  wire n616_o;
  wire n617_o;
  wire [1:0] n618_o;
  reg n620_o;
  wire [3:0] n627_o;
  wire [3:0] n628_o;
  wire [3:0] n629_o;
  wire n637_o;
  wire n639_o;
  wire n640_o;
  wire n642_o;
  wire n643_o;
  wire n645_o;
  wire n646_o;
  wire n648_o;
  wire n649_o;
  wire n651_o;
  wire n652_o;
  reg n655_o;
  wire [7:0] n658_o;
  wire [7:0] n660_o;
  reg [7:0] n661_q;
  wire [7:0] n662_o;
  reg [7:0] n663_q;
  wire [7:0] n664_o;
  reg [7:0] n665_q;
  wire [7:0] n666_o;
  assign data_o = n658_o;
  assign carry_o = n496_o;
  assign aux_carry_o = n620_o;
  assign da_overflow_o = n655_o;
  /* alu.vhd:99:10  */
  assign accumulator_q = n661_q; // (signal)
  /* alu.vhd:100:10  */
  assign accu_shadow_q = n663_q; // (signal)
  /* alu.vhd:101:10  */
  assign temp_req_q = n665_q; // (signal)
  /* alu.vhd:103:10  */
  assign in_a_s = accu_shadow_q; // (signal)
  /* alu.vhd:104:10  */
  assign in_b_s = temp_req_q; // (signal)
  /* alu.vhd:106:10  */
  assign data_s = n666_o; // (signal)
  /* alu.vhd:108:10  */
  assign add_result_s = n595_o; // (signal)
  /* alu.vhd:122:14  */
  assign n417_o = ~res_i;
  /* alu.vhd:132:52  */
  assign n419_o = data_i[3:0];
  /* t48_core.vhd:568:26  */
  assign n420_o = data_i[3:0];
  /* alu.vhd:131:11  */
  assign n421_o = accu_low_i ? n419_o : n420_o;
  /* t48_core.vhd:551:5  */
  assign n422_o = data_i[7:4];
  /* t48_core.vhd:551:5  */
  assign n423_o = accumulator_q[7:4];
  /* alu.vhd:131:11  */
  assign n424_o = accu_low_i ? n423_o : n422_o;
  /* t48_core.vhd:551:5  */
  assign n425_o = {n424_o, n421_o};
  /* alu.vhd:138:9  */
  assign n427_o = write_shadow_i ? data_i : accumulator_q;
  /* alu.vhd:152:9  */
  assign n428_o = write_temp_reg_i ? data_i : temp_req_q;
  /* alu.vhd:149:9  */
  assign n430_o = p60_temp_reg_i ? 8'b01100000 : n428_o;
  /* alu.vhd:146:9  */
  assign n432_o = p06_temp_reg_i ? 8'b00000110 : n430_o;
  /* alu.vhd:128:7  */
  assign n433_o = en_clk_i & write_accu_i;
  /* alu.vhd:203:26  */
  assign n447_o = in_a_s & in_b_s;
  /* alu.vhd:202:7  */
  assign n449_o = alu_op_i == 4'b0000;
  /* alu.vhd:207:26  */
  assign n450_o = in_a_s | in_b_s;
  /* alu.vhd:206:7  */
  assign n452_o = alu_op_i == 4'b0001;
  /* alu.vhd:211:26  */
  assign n453_o = in_a_s ^ in_b_s;
  /* alu.vhd:210:7  */
  assign n455_o = alu_op_i == 4'b0010;
  /* alu.vhd:215:32  */
  assign n456_o = add_result_s[7:0];
  /* alu.vhd:216:32  */
  assign n457_o = add_result_s[8];
  /* alu.vhd:214:7  */
  assign n459_o = alu_op_i == 4'b1010;
  /* alu.vhd:220:19  */
  assign n460_o = ~in_a_s;
  /* alu.vhd:219:7  */
  assign n462_o = alu_op_i == 4'b0011;
  /* alu.vhd:223:7  */
  assign n464_o = alu_op_i == 4'b0100;
  /* alu.vhd:228:37  */
  assign n465_o = in_a_s[6:0];
  /* alu.vhd:229:37  */
  assign n466_o = in_a_s[7];
  /* alu.vhd:234:37  */
  assign n467_o = in_a_s[7];
  /* alu.vhd:231:9  */
  assign n468_o = use_carry_i ? carry_i : n467_o;
  /* alu.vhd:227:7  */
  assign n470_o = alu_op_i == 4'b0101;
  /* alu.vhd:239:37  */
  assign n471_o = in_a_s[7:1];
  /* alu.vhd:240:37  */
  assign n472_o = in_a_s[0];
  /* alu.vhd:245:37  */
  assign n473_o = in_a_s[0];
  /* alu.vhd:242:9  */
  assign n474_o = use_carry_i ? carry_i : n473_o;
  /* alu.vhd:238:7  */
  assign n476_o = alu_op_i == 4'b0110;
  /* alu.vhd:250:37  */
  assign n477_o = in_a_s[7:4];
  /* alu.vhd:251:37  */
  assign n478_o = in_a_s[3:0];
  /* alu.vhd:249:7  */
  assign n480_o = alu_op_i == 4'b0111;
  /* alu.vhd:255:31  */
  assign n481_o = add_result_s[7:0];
  /* alu.vhd:254:7  */
  assign n483_o = alu_op_i == 4'b1000;
  /* alu.vhd:259:31  */
  assign n484_o = add_result_s[7:0];
  /* alu.vhd:258:7  */
  assign n486_o = alu_op_i == 4'b1001;
  /* alu.vhd:263:25  */
  assign n487_o = in_b_s[7:4];
  /* alu.vhd:263:46  */
  assign n488_o = in_a_s[3:0];
  /* alu.vhd:263:38  */
  assign n489_o = {n487_o, n488_o};
  /* alu.vhd:262:7  */
  assign n491_o = alu_op_i == 4'b1011;
  /* alu.vhd:266:7  */
  assign n493_o = alu_op_i == 4'b1100;
  /* t48_core.vhd:418:33  */
  assign n494_o = {n493_o, n491_o, n486_o, n483_o, n480_o, n476_o, n470_o, n464_o, n462_o, n459_o, n455_o, n452_o, n449_o};
  /* alu.vhd:200:5  */
  always @*
    case (n494_o)
      13'b1000000000000: n496_o = 1'b0;
      13'b0100000000000: n496_o = 1'b0;
      13'b0010000000000: n496_o = 1'b0;
      13'b0001000000000: n496_o = 1'b0;
      13'b0000100000000: n496_o = 1'b0;
      13'b0000010000000: n496_o = n472_o;
      13'b0000001000000: n496_o = n466_o;
      13'b0000000100000: n496_o = 1'b0;
      13'b0000000010000: n496_o = 1'b0;
      13'b0000000001000: n496_o = n457_o;
      13'b0000000000100: n496_o = 1'b0;
      13'b0000000000010: n496_o = 1'b0;
      13'b0000000000001: n496_o = 1'b0;
      default: n496_o = 1'b0;
    endcase
  /* t48_core.vhd:414:33  */
  assign n498_o = n447_o[0];
  /* t48_core.vhd:413:33  */
  assign n499_o = n450_o[0];
  /* t48_core.vhd:412:33  */
  assign n500_o = n453_o[0];
  /* t48_core.vhd:411:33  */
  assign n501_o = n456_o[0];
  /* t48_core.vhd:410:33  */
  assign n502_o = n460_o[0];
  /* t48_core.vhd:408:33  */
  assign n504_o = n471_o[0];
  /* t48_core.vhd:407:33  */
  assign n505_o = n477_o[0];
  /* t48_core.vhd:405:33  */
  assign n506_o = n481_o[0];
  /* t48_core.vhd:392:3  */
  assign n507_o = n484_o[0];
  /* t48_core.vhd:392:3  */
  assign n508_o = n489_o[0];
  /* t48_core.vhd:392:3  */
  assign n509_o = in_a_s[0];
  /* alu.vhd:200:5  */
  always @*
    case (n494_o)
      13'b1000000000000: n511_o = n509_o;
      13'b0100000000000: n511_o = n508_o;
      13'b0010000000000: n511_o = n507_o;
      13'b0001000000000: n511_o = n506_o;
      13'b0000100000000: n511_o = n505_o;
      13'b0000010000000: n511_o = n504_o;
      13'b0000001000000: n511_o = n468_o;
      13'b0000000100000: n511_o = 1'b0;
      13'b0000000010000: n511_o = n502_o;
      13'b0000000001000: n511_o = n501_o;
      13'b0000000000100: n511_o = n500_o;
      13'b0000000000010: n511_o = n499_o;
      13'b0000000000001: n511_o = n498_o;
      default: n511_o = 1'b0;
    endcase
  /* t48_core.vhd:392:3  */
  assign n512_o = n447_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n513_o = n450_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n514_o = n453_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n515_o = n456_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n516_o = n460_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n518_o = n465_o[2:0];
  /* t48_core.vhd:392:3  */
  assign n519_o = n471_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n520_o = n477_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n521_o = n481_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n522_o = n484_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n523_o = n489_o[3:1];
  /* t48_core.vhd:392:3  */
  assign n524_o = in_a_s[3:1];
  /* alu.vhd:200:5  */
  always @*
    case (n494_o)
      13'b1000000000000: n526_o = n524_o;
      13'b0100000000000: n526_o = n523_o;
      13'b0010000000000: n526_o = n522_o;
      13'b0001000000000: n526_o = n521_o;
      13'b0000100000000: n526_o = n520_o;
      13'b0000010000000: n526_o = n519_o;
      13'b0000001000000: n526_o = n518_o;
      13'b0000000100000: n526_o = 3'b000;
      13'b0000000010000: n526_o = n516_o;
      13'b0000000001000: n526_o = n515_o;
      13'b0000000000100: n526_o = n514_o;
      13'b0000000000010: n526_o = n513_o;
      13'b0000000000001: n526_o = n512_o;
      default: n526_o = 3'b000;
    endcase
  /* t48_core.vhd:392:3  */
  assign n527_o = n447_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n528_o = n450_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n529_o = n453_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n530_o = n456_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n531_o = n460_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n533_o = n465_o[5:3];
  /* t48_core.vhd:392:3  */
  assign n534_o = n471_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n535_o = n478_o[2:0];
  /* t48_core.vhd:392:3  */
  assign n536_o = n481_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n537_o = n484_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n538_o = n489_o[6:4];
  /* t48_core.vhd:392:3  */
  assign n539_o = in_a_s[6:4];
  /* alu.vhd:200:5  */
  always @*
    case (n494_o)
      13'b1000000000000: n541_o = n539_o;
      13'b0100000000000: n541_o = n538_o;
      13'b0010000000000: n541_o = n537_o;
      13'b0001000000000: n541_o = n536_o;
      13'b0000100000000: n541_o = n535_o;
      13'b0000010000000: n541_o = n534_o;
      13'b0000001000000: n541_o = n533_o;
      13'b0000000100000: n541_o = 3'b000;
      13'b0000000010000: n541_o = n531_o;
      13'b0000000001000: n541_o = n530_o;
      13'b0000000000100: n541_o = n529_o;
      13'b0000000000010: n541_o = n528_o;
      13'b0000000000001: n541_o = n527_o;
      default: n541_o = 3'b000;
    endcase
  /* t48_core.vhd:392:3  */
  assign n542_o = n447_o[7];
  /* t48_core.vhd:392:3  */
  assign n543_o = n450_o[7];
  /* t48_core.vhd:392:3  */
  assign n544_o = n453_o[7];
  /* t48_core.vhd:392:3  */
  assign n545_o = n456_o[7];
  /* t48_core.vhd:392:3  */
  assign n546_o = n460_o[7];
  /* t48_core.vhd:392:3  */
  assign n548_o = n465_o[6];
  /* t48_core.vhd:392:3  */
  assign n549_o = n478_o[3];
  /* t48_core.vhd:392:3  */
  assign n550_o = n481_o[7];
  /* t48_core.vhd:392:3  */
  assign n551_o = n484_o[7];
  /* t48_core.vhd:392:3  */
  assign n552_o = n489_o[7];
  /* t48_core.vhd:392:3  */
  assign n553_o = in_a_s[7];
  /* alu.vhd:200:5  */
  always @*
    case (n494_o)
      13'b1000000000000: n555_o = n553_o;
      13'b0100000000000: n555_o = n552_o;
      13'b0010000000000: n555_o = n551_o;
      13'b0001000000000: n555_o = n550_o;
      13'b0000100000000: n555_o = n549_o;
      13'b0000010000000: n555_o = n474_o;
      13'b0000001000000: n555_o = n548_o;
      13'b0000000100000: n555_o = 1'b0;
      13'b0000000010000: n555_o = n546_o;
      13'b0000000001000: n555_o = n545_o;
      13'b0000000000100: n555_o = n544_o;
      13'b0000000000010: n555_o = n543_o;
      13'b0000000000001: n555_o = n542_o;
      default: n555_o = 1'b0;
    endcase
  /* alu.vhd:307:20  */
  assign n567_o = carry_i & use_carry_i;
  /* alu.vhd:307:5  */
  assign n570_o = n567_o ? 1'b1 : 1'b0;
  /* t48_core.vhd:347:3  */
  assign n572_o = n571_o[8:1];
  /* alu.vhd:313:20  */
  assign n574_o = {1'b0, in_a_s};
  /* alu.vhd:314:20  */
  assign n576_o = {1'b0, in_b_s};
  /* t48_core.vhd:338:25  */
  assign n579_o = n578_o[8:1];
  /* alu.vhd:317:7  */
  assign n581_o = alu_op_i == 4'b1001;
  /* alu.vhd:320:7  */
  assign n583_o = alu_op_i == 4'b1000;
  /* t48_core.vhd:321:3  */
  assign n584_o = {n583_o, n581_o};
  /* t48_core.vhd:321:3  */
  assign n586_o = n576_o[0];
  /* alu.vhd:316:5  */
  always @*
    case (n584_o)
      2'b10: n587_o = 1'b1;
      2'b01: n587_o = 1'b1;
      default: n587_o = n586_o;
    endcase
  /* t48_core.vhd:321:3  */
  assign n589_o = n576_o[8:1];
  /* alu.vhd:316:5  */
  always @*
    case (n584_o)
      2'b10: n590_o = 8'b11111111;
      2'b01: n590_o = n579_o;
      default: n590_o = n589_o;
    endcase
  /* t48_core.vhd:307:3  */
  assign n592_o = {n590_o, n587_o};
  /* alu.vhd:327:35  */
  assign n593_o = n574_o + n592_o;
  /* t48_core.vhd:297:29  */
  assign n594_o = {n572_o, n570_o};
  /* alu.vhd:328:35  */
  assign n595_o = n593_o + n594_o;
  /* alu.vhd:334:32  */
  assign n596_o = in_a_s[4];
  /* alu.vhd:334:44  */
  assign n597_o = in_b_s[4];
  /* alu.vhd:334:36  */
  assign n598_o = {n596_o, n597_o};
  /* alu.vhd:339:20  */
  assign n599_o = n595_o[4];
  /* alu.vhd:339:9  */
  assign n602_o = n599_o ? 1'b1 : 1'b0;
  /* alu.vhd:338:7  */
  assign n604_o = n598_o == 2'b00;
  /* alu.vhd:338:17  */
  assign n606_o = n598_o == 2'b11;
  /* alu.vhd:338:17  */
  assign n607_o = n604_o | n606_o;
  /* alu.vhd:344:20  */
  assign n608_o = n595_o[4];
  /* alu.vhd:344:24  */
  assign n609_o = ~n608_o;
  /* alu.vhd:344:9  */
  assign n612_o = n609_o ? 1'b1 : 1'b0;
  /* alu.vhd:343:7  */
  assign n614_o = n598_o == 2'b01;
  /* alu.vhd:343:17  */
  assign n616_o = n598_o == 2'b10;
  /* alu.vhd:343:17  */
  assign n617_o = n614_o | n616_o;
  /* t48_core.vhd:87:5  */
  assign n618_o = {n617_o, n607_o};
  /* alu.vhd:337:5  */
  always @*
    case (n618_o)
      2'b10: n620_o = n612_o;
      2'b01: n620_o = n602_o;
      default: n620_o = 1'b0;
    endcase
  /* alu.vhd:389:35  */
  assign n627_o = accu_shadow_q[7:4];
  /* alu.vhd:391:35  */
  assign n628_o = accu_shadow_q[3:0];
  /* alu.vhd:388:5  */
  assign n629_o = da_high_i ? n627_o : n628_o;
  /* alu.vhd:373:9  */
  assign n637_o = n629_o == 4'b1010;
  /* alu.vhd:373:21  */
  assign n639_o = n629_o == 4'b1011;
  /* alu.vhd:373:21  */
  assign n640_o = n637_o | n639_o;
  /* alu.vhd:374:21  */
  assign n642_o = n629_o == 4'b1100;
  /* alu.vhd:374:21  */
  assign n643_o = n640_o | n642_o;
  /* alu.vhd:375:21  */
  assign n645_o = n629_o == 4'b1101;
  /* alu.vhd:375:21  */
  assign n646_o = n643_o | n645_o;
  /* alu.vhd:376:21  */
  assign n648_o = n629_o == 4'b1110;
  /* alu.vhd:376:21  */
  assign n649_o = n646_o | n648_o;
  /* alu.vhd:377:21  */
  assign n651_o = n629_o == 4'b1111;
  /* alu.vhd:377:21  */
  assign n652_o = n649_o | n651_o;
  /* alu.vhd:372:7  */
  always @*
    case (n652_o)
      1'b1: n655_o = 1'b1;
      default: n655_o = 1'b0;
    endcase
  /* alu.vhd:412:13  */
  assign n658_o = read_alu_i ? data_s : 8'b11111111;
  /* alu.vhd:127:5  */
  assign n660_o = n433_o ? n425_o : accumulator_q;
  /* alu.vhd:127:5  */
  always @(posedge clk_i or posedge n417_o)
    if (n417_o)
      n661_q <= 8'b00000000;
    else
      n661_q <= n660_o;
  /* alu.vhd:127:5  */
  assign n662_o = en_clk_i ? n427_o : accu_shadow_q;
  /* alu.vhd:127:5  */
  always @(posedge clk_i or posedge n417_o)
    if (n417_o)
      n663_q <= 8'b00000000;
    else
      n663_q <= n662_o;
  /* alu.vhd:127:5  */
  assign n664_o = en_clk_i ? n432_o : temp_req_q;
  /* alu.vhd:127:5  */
  always @(posedge clk_i or posedge n417_o)
    if (n417_o)
      n665_q <= 8'b00000000;
    else
      n665_q <= n664_o;
  /* alu.vhd:122:5  */
  assign n666_o = {n555_o, n541_o, n526_o, n511_o};
endmodule

module t48_core
  (input  xtal_i,
   input  xtal_en_i,
   input  reset_i,
   input  t0_i,
   input  int_n_i,
   input  ea_i,
   input  [7:0] db_i,
   input  t1_i,
   input  [7:0] p2_i,
   input  [7:0] p1_i,
   input  clk_i,
   input  en_clk_i,
   input  [7:0] dmem_data_i,
   input  [7:0] pmem_data_i,
   output t0_o,
   output t0_dir_o,
   output rd_n_o,
   output psen_n_o,
   output wr_n_o,
   output ale_o,
   output [7:0] db_o,
   output db_dir_o,
   output [7:0] p2_o,
   output p2l_low_imp_o,
   output p2h_low_imp_o,
   output [7:0] p1_o,
   output p1_low_imp_o,
   output prog_n_o,
   output xtal3_o,
   output [7:0] dmem_addr_o,
   output dmem_we_o,
   output [7:0] dmem_data_o,
   output [11:0] pmem_addr_o);
  wire [7:0] t48_data_s;
  wire xtal_en_s;
  wire en_clk_s;
  wire t0_s;
  wire t1_s;
  wire [7:0] alu_data_s;
  wire alu_write_accu_s;
  wire alu_write_shadow_s;
  wire alu_write_temp_reg_s;
  wire alu_read_alu_s;
  wire alu_carry_s;
  wire alu_aux_carry_s;
  wire [3:0] alu_op_s;
  wire alu_use_carry_s;
  wire alu_da_high_s;
  wire alu_da_overflow_s;
  wire alu_accu_low_s;
  wire alu_p06_temp_reg_s;
  wire alu_p60_temp_reg_s;
  wire bus_write_bus_s;
  wire bus_read_bus_s;
  wire bus_output_pcl_s;
  wire bus_bidir_bus_s;
  wire [7:0] bus_data_s;
  wire clk_multi_cycle_s;
  wire clk_assert_psen_s;
  wire clk_assert_prog_s;
  wire clk_assert_rd_s;
  wire clk_assert_wr_s;
  wire [2:0] clk_mstate_s;
  wire clk_second_cycle_s;
  wire psen_s;
  wire prog_s;
  wire rd_s;
  wire wr_s;
  wire ale_s;
  wire xtal3_s;
  wire cnd_compute_take_s;
  wire [3:0] cnd_branch_cond_s;
  wire cnd_take_branch_s;
  wire [2:0] cnd_comp_value_s;
  wire cnd_f1_s;
  wire cnd_tf_s;
  wire dm_write_dmem_addr_s;
  wire dm_write_dmem_s;
  wire dm_read_dmem_s;
  wire [1:0] dm_addr_type_s;
  wire [7:0] dm_data_s;
  wire [7:0] dec_data_s;
  wire p1_write_p1_s;
  wire p1_read_p1_s;
  wire p1_read_reg_s;
  wire [7:0] p1_data_s;
  wire p2_write_p2_s;
  wire p2_write_exp_s;
  wire p2_read_p2_s;
  wire p2_read_reg_s;
  wire p2_read_exp_s;
  wire p2_output_pch_s;
  wire [7:0] p2_data_s;
  wire pm_write_pcl_s;
  wire pm_read_pcl_s;
  wire pm_write_pch_s;
  wire pm_read_pch_s;
  wire pm_read_pmem_s;
  wire pm_inc_pc_s;
  wire pm_write_pmem_addr_s;
  wire [7:0] pm_data_s;
  wire [1:0] pm_addr_type_s;
  wire [11:0] pmem_addr_s;
  wire psw_read_psw_s;
  wire psw_read_sp_s;
  wire psw_write_psw_s;
  wire psw_write_sp_s;
  wire psw_carry_s;
  wire psw_aux_carry_s;
  wire psw_f0_s;
  wire psw_bs_s;
  wire psw_special_data_s;
  wire psw_inc_stackp_s;
  wire psw_dec_stackp_s;
  wire psw_write_carry_s;
  wire psw_write_aux_carry_s;
  wire psw_write_f0_s;
  wire psw_write_bs_s;
  wire [7:0] psw_data_s;
  wire tim_overflow_s;
  wire tim_of_s;
  wire tim_read_timer_s;
  wire tim_write_timer_s;
  wire tim_start_t_s;
  wire tim_start_cnt_s;
  wire tim_stop_tcnt_s;
  wire [7:0] tim_data_s;
  wire n26_o;
  wire n34_o;
  wire [7:0] alu_b_n35;
  wire alu_b_n36;
  wire alu_b_n37;
  wire alu_b_n38;
  wire [7:0] alu_b_data_o;
  wire alu_b_carry_o;
  wire alu_b_aux_carry_o;
  wire alu_b_da_overflow_o;
  wire [7:0] bus_mux_b_n47;
  wire [7:0] bus_mux_b_data_o;
  wire clock_ctrl_b_n50;
  wire clock_ctrl_b_n51;
  wire [2:0] clock_ctrl_b_n52;
  wire clock_ctrl_b_n53;
  wire clock_ctrl_b_n54;
  wire clock_ctrl_b_n55;
  wire clock_ctrl_b_n56;
  wire clock_ctrl_b_n57;
  wire clock_ctrl_b_n58;
  wire clock_ctrl_b_xtal3_o;
  wire clock_ctrl_b_t0_o;
  wire [2:0] clock_ctrl_b_mstate_o;
  wire clock_ctrl_b_second_cycle_o;
  wire clock_ctrl_b_ale_o;
  wire clock_ctrl_b_psen_o;
  wire clock_ctrl_b_prog_o;
  wire clock_ctrl_b_rd_o;
  wire clock_ctrl_b_wr_o;
  wire cond_branch_b_n77;
  localparam n78_o = 1'b0;
  localparam n79_o = 1'b0;
  wire cond_branch_b_take_branch_o;
  wire [7:0] use_db_bus_db_bus_b_n82;
  wire [7:0] n83_o;
  wire [7:0] use_db_bus_db_bus_b_n84;
  wire use_db_bus_db_bus_b_n85;
  wire [7:0] use_db_bus_db_bus_b_data_o;
  wire [7:0] use_db_bus_db_bus_b_db_o;
  wire use_db_bus_db_bus_b_db_dir_o;
  wire decoder_b_n92;
  wire [7:0] decoder_b_n93;
  wire decoder_b_n94;
  wire decoder_b_n95;
  wire decoder_b_n96;
  wire decoder_b_n97;
  wire decoder_b_n98;
  wire decoder_b_n99;
  localparam n100_o = 1'b0;
  localparam n101_o = 1'b0;
  wire decoder_b_n106;
  wire decoder_b_n107;
  wire decoder_b_n108;
  wire decoder_b_n109;
  wire decoder_b_n110;
  wire decoder_b_n111;
  wire decoder_b_n112;
  wire decoder_b_n113;
  wire decoder_b_n114;
  wire decoder_b_n115;
  wire decoder_b_n116;
  wire decoder_b_n117;
  wire decoder_b_n118;
  wire decoder_b_n119;
  wire decoder_b_n120;
  wire decoder_b_n121;
  wire decoder_b_n122;
  wire [3:0] decoder_b_n123;
  wire decoder_b_n124;
  wire decoder_b_n125;
  wire decoder_b_n126;
  wire decoder_b_n127;
  wire decoder_b_n128;
  wire decoder_b_n129;
  wire decoder_b_n130;
  wire decoder_b_n131;
  wire decoder_b_n132;
  wire decoder_b_n133;
  wire decoder_b_n134;
  wire decoder_b_n135;
  wire decoder_b_n136;
  wire [3:0] decoder_b_n137;
  wire [2:0] decoder_b_n138;
  wire decoder_b_n139;
  wire decoder_b_n140;
  wire [1:0] decoder_b_n141;
  wire decoder_b_n142;
  wire decoder_b_n143;
  wire decoder_b_n144;
  wire decoder_b_n145;
  wire decoder_b_n146;
  wire decoder_b_n147;
  wire decoder_b_n148;
  wire decoder_b_n149;
  wire decoder_b_n150;
  wire decoder_b_n151;
  wire decoder_b_n152;
  wire [1:0] decoder_b_n153;
  wire decoder_b_n154;
  wire decoder_b_n155;
  wire decoder_b_n156;
  wire decoder_b_n157;
  wire decoder_b_n158;
  wire decoder_b_n159;
  wire decoder_b_n160;
  wire decoder_b_t0_dir_o;
  wire [7:0] decoder_b_data_o;
  wire decoder_b_alu_write_accu_o;
  wire decoder_b_alu_write_shadow_o;
  wire decoder_b_alu_write_temp_reg_o;
  wire decoder_b_alu_read_alu_o;
  wire decoder_b_bus_write_bus_o;
  wire decoder_b_bus_read_bus_o;
  wire decoder_b_bus_ibf_int_o;
  wire decoder_b_bus_en_dma_o;
  wire decoder_b_bus_en_flags_o;
  wire decoder_b_bus_write_sts_o;
  wire decoder_b_dm_write_dmem_addr_o;
  wire decoder_b_dm_write_dmem_o;
  wire decoder_b_dm_read_dmem_o;
  wire decoder_b_p1_write_p1_o;
  wire decoder_b_p1_read_p1_o;
  wire decoder_b_p2_write_p2_o;
  wire decoder_b_p2_write_exp_o;
  wire decoder_b_p2_read_p2_o;
  wire decoder_b_p2_read_exp_o;
  wire decoder_b_pm_write_pcl_o;
  wire decoder_b_pm_read_pcl_o;
  wire decoder_b_pm_write_pch_o;
  wire decoder_b_pm_read_pch_o;
  wire decoder_b_pm_read_pmem_o;
  wire decoder_b_psw_read_psw_o;
  wire decoder_b_psw_read_sp_o;
  wire decoder_b_psw_write_psw_o;
  wire decoder_b_psw_write_sp_o;
  wire [3:0] decoder_b_alu_op_o;
  wire decoder_b_alu_use_carry_o;
  wire decoder_b_alu_da_high_o;
  wire decoder_b_alu_accu_low_o;
  wire decoder_b_alu_p06_temp_reg_o;
  wire decoder_b_alu_p60_temp_reg_o;
  wire decoder_b_bus_output_pcl_o;
  wire decoder_b_bus_bidir_bus_o;
  wire decoder_b_clk_multi_cycle_o;
  wire decoder_b_clk_assert_psen_o;
  wire decoder_b_clk_assert_prog_o;
  wire decoder_b_clk_assert_rd_o;
  wire decoder_b_clk_assert_wr_o;
  wire decoder_b_cnd_compute_take_o;
  wire [3:0] decoder_b_cnd_branch_cond_o;
  wire [2:0] decoder_b_cnd_comp_value_o;
  wire decoder_b_cnd_f1_o;
  wire decoder_b_cnd_tf_o;
  wire [1:0] decoder_b_dm_addr_type_o;
  wire decoder_b_p1_read_reg_o;
  wire decoder_b_p2_read_reg_o;
  wire decoder_b_p2_output_pch_o;
  wire decoder_b_pm_inc_pc_o;
  wire decoder_b_pm_write_pmem_addr_o;
  wire [1:0] decoder_b_pm_addr_type_o;
  wire decoder_b_psw_special_data_o;
  wire decoder_b_psw_inc_stackp_o;
  wire decoder_b_psw_dec_stackp_o;
  wire decoder_b_psw_write_carry_o;
  wire decoder_b_psw_write_aux_carry_o;
  wire decoder_b_psw_write_f0_o;
  wire decoder_b_psw_write_bs_o;
  wire decoder_b_tim_read_timer_o;
  wire decoder_b_tim_write_timer_o;
  wire decoder_b_tim_start_t_o;
  wire decoder_b_tim_start_cnt_o;
  wire decoder_b_tim_stop_tcnt_o;
  wire [7:0] dmem_ctrl_b_n291;
  wire [7:0] dmem_ctrl_b_n292;
  wire dmem_ctrl_b_n293;
  wire [7:0] dmem_ctrl_b_n294;
  wire [7:0] dmem_ctrl_b_data_o;
  wire [7:0] dmem_ctrl_b_dmem_addr_o;
  wire dmem_ctrl_b_dmem_we_o;
  wire [7:0] dmem_ctrl_b_dmem_data_o;
  wire [7:0] use_timer_timer_b_n303;
  wire use_timer_timer_b_n304;
  wire [7:0] use_timer_timer_b_data_o;
  wire use_timer_timer_b_overflow_o;
  wire n316_o;
  wire [7:0] use_p1_p1_b_n317;
  wire [7:0] use_p1_p1_b_n318;
  wire use_p1_p1_b_n319;
  wire [7:0] use_p1_p1_b_data_o;
  wire [7:0] use_p1_p1_b_p1_o;
  wire use_p1_p1_b_p1_low_imp_o;
  wire [7:0] use_p2_p2_b_n326;
  wire [3:0] n327_o;
  wire [7:0] use_p2_p2_b_n328;
  wire use_p2_p2_b_n329;
  wire use_p2_p2_b_n330;
  wire [7:0] use_p2_p2_b_data_o;
  wire [7:0] use_p2_p2_b_p2_o;
  wire use_p2_p2_b_p2l_low_imp_o;
  wire use_p2_p2_b_p2h_low_imp_o;
  wire [7:0] pmem_ctrl_b_n339;
  wire [11:0] pmem_ctrl_b_n340;
  wire [7:0] pmem_ctrl_b_data_o;
  wire [11:0] pmem_ctrl_b_pmem_addr_o;
  wire [7:0] psw_b_n345;
  wire psw_b_n346;
  wire psw_b_n347;
  wire psw_b_n348;
  wire psw_b_n349;
  wire [7:0] psw_b_data_o;
  wire psw_b_carry_o;
  wire psw_b_aux_carry_o;
  wire psw_b_f0_o;
  wire psw_b_bs_o;
  wire n367_o;
  wire n369_o;
  wire n376_o;
  wire n378_o;
  wire n385_o;
  wire n387_o;
  wire n394_o;
  wire n396_o;
  wire n403_o;
  wire n411_o;
  assign t0_o = clock_ctrl_b_n51;
  assign t0_dir_o = decoder_b_n92;
  assign rd_n_o = n394_o;
  assign psen_n_o = n376_o;
  assign wr_n_o = n403_o;
  assign ale_o = n367_o;
  assign db_o = use_db_bus_db_bus_b_n84;
  assign db_dir_o = use_db_bus_db_bus_b_n85;
  assign p2_o = use_p2_p2_b_n328;
  assign p2l_low_imp_o = use_p2_p2_b_n329;
  assign p2h_low_imp_o = use_p2_p2_b_n330;
  assign p1_o = use_p1_p1_b_n318;
  assign p1_low_imp_o = use_p1_p1_b_n319;
  assign prog_n_o = n385_o;
  assign xtal3_o = n411_o;
  assign dmem_addr_o = dmem_ctrl_b_n292;
  assign dmem_we_o = dmem_ctrl_b_n293;
  assign dmem_data_o = dmem_ctrl_b_n294;
  assign pmem_addr_o = pmem_addr_s;
  /* t48_core.vhd:136:10  */
  assign t48_data_s = bus_mux_b_n47; // (signal)
  /* t48_core.vhd:138:10  */
  assign xtal_en_s = n26_o; // (signal)
  /* t48_core.vhd:139:10  */
  assign en_clk_s = n34_o; // (signal)
  /* t48_core.vhd:141:10  */
  assign t0_s = t0_i; // (signal)
  /* t48_core.vhd:141:16  */
  assign t1_s = t1_i; // (signal)
  /* t48_core.vhd:144:10  */
  assign alu_data_s = alu_b_n35; // (signal)
  /* t48_core.vhd:145:10  */
  assign alu_write_accu_s = decoder_b_n94; // (signal)
  /* t48_core.vhd:146:10  */
  assign alu_write_shadow_s = decoder_b_n95; // (signal)
  /* t48_core.vhd:147:10  */
  assign alu_write_temp_reg_s = decoder_b_n96; // (signal)
  /* t48_core.vhd:148:10  */
  assign alu_read_alu_s = decoder_b_n97; // (signal)
  /* t48_core.vhd:149:10  */
  assign alu_carry_s = alu_b_n36; // (signal)
  /* t48_core.vhd:150:10  */
  assign alu_aux_carry_s = alu_b_n37; // (signal)
  /* t48_core.vhd:151:10  */
  assign alu_op_s = decoder_b_n123; // (signal)
  /* t48_core.vhd:152:10  */
  assign alu_use_carry_s = decoder_b_n128; // (signal)
  /* t48_core.vhd:153:10  */
  assign alu_da_high_s = decoder_b_n124; // (signal)
  /* t48_core.vhd:154:10  */
  assign alu_da_overflow_s = alu_b_n38; // (signal)
  /* t48_core.vhd:155:10  */
  assign alu_accu_low_s = decoder_b_n125; // (signal)
  /* t48_core.vhd:156:10  */
  assign alu_p06_temp_reg_s = decoder_b_n126; // (signal)
  /* t48_core.vhd:157:10  */
  assign alu_p60_temp_reg_s = decoder_b_n127; // (signal)
  /* t48_core.vhd:160:10  */
  assign bus_write_bus_s = decoder_b_n98; // (signal)
  /* t48_core.vhd:161:10  */
  assign bus_read_bus_s = decoder_b_n99; // (signal)
  /* t48_core.vhd:162:10  */
  assign bus_output_pcl_s = decoder_b_n129; // (signal)
  /* t48_core.vhd:163:10  */
  assign bus_bidir_bus_s = decoder_b_n130; // (signal)
  /* t48_core.vhd:164:10  */
  assign bus_data_s = use_db_bus_db_bus_b_n82; // (signal)
  /* t48_core.vhd:167:10  */
  assign clk_multi_cycle_s = decoder_b_n131; // (signal)
  /* t48_core.vhd:168:10  */
  assign clk_assert_psen_s = decoder_b_n132; // (signal)
  /* t48_core.vhd:169:10  */
  assign clk_assert_prog_s = decoder_b_n133; // (signal)
  /* t48_core.vhd:170:10  */
  assign clk_assert_rd_s = decoder_b_n134; // (signal)
  /* t48_core.vhd:171:10  */
  assign clk_assert_wr_s = decoder_b_n135; // (signal)
  /* t48_core.vhd:172:10  */
  assign clk_mstate_s = clock_ctrl_b_n52; // (signal)
  /* t48_core.vhd:173:10  */
  assign clk_second_cycle_s = clock_ctrl_b_n53; // (signal)
  /* t48_core.vhd:174:10  */
  assign psen_s = clock_ctrl_b_n55; // (signal)
  /* t48_core.vhd:175:10  */
  assign prog_s = clock_ctrl_b_n56; // (signal)
  /* t48_core.vhd:176:10  */
  assign rd_s = clock_ctrl_b_n57; // (signal)
  /* t48_core.vhd:177:10  */
  assign wr_s = clock_ctrl_b_n58; // (signal)
  /* t48_core.vhd:178:10  */
  assign ale_s = clock_ctrl_b_n54; // (signal)
  /* t48_core.vhd:179:10  */
  assign xtal3_s = clock_ctrl_b_n50; // (signal)
  /* t48_core.vhd:182:10  */
  assign cnd_compute_take_s = decoder_b_n136; // (signal)
  /* t48_core.vhd:183:10  */
  assign cnd_branch_cond_s = decoder_b_n137; // (signal)
  /* t48_core.vhd:184:10  */
  assign cnd_take_branch_s = cond_branch_b_n77; // (signal)
  /* t48_core.vhd:185:10  */
  assign cnd_comp_value_s = decoder_b_n138; // (signal)
  /* t48_core.vhd:186:10  */
  assign cnd_f1_s = decoder_b_n139; // (signal)
  /* t48_core.vhd:187:10  */
  assign cnd_tf_s = decoder_b_n140; // (signal)
  /* t48_core.vhd:190:10  */
  assign dm_write_dmem_addr_s = decoder_b_n106; // (signal)
  /* t48_core.vhd:191:10  */
  assign dm_write_dmem_s = decoder_b_n107; // (signal)
  /* t48_core.vhd:192:10  */
  assign dm_read_dmem_s = decoder_b_n108; // (signal)
  /* t48_core.vhd:193:10  */
  assign dm_addr_type_s = decoder_b_n141; // (signal)
  /* t48_core.vhd:194:10  */
  assign dm_data_s = dmem_ctrl_b_n291; // (signal)
  /* t48_core.vhd:197:10  */
  assign dec_data_s = decoder_b_n93; // (signal)
  /* t48_core.vhd:200:10  */
  assign p1_write_p1_s = decoder_b_n109; // (signal)
  /* t48_core.vhd:201:10  */
  assign p1_read_p1_s = decoder_b_n110; // (signal)
  /* t48_core.vhd:202:10  */
  assign p1_read_reg_s = decoder_b_n147; // (signal)
  /* t48_core.vhd:203:10  */
  assign p1_data_s = use_p1_p1_b_n317; // (signal)
  /* t48_core.vhd:206:10  */
  assign p2_write_p2_s = decoder_b_n111; // (signal)
  /* t48_core.vhd:207:10  */
  assign p2_write_exp_s = decoder_b_n112; // (signal)
  /* t48_core.vhd:208:10  */
  assign p2_read_p2_s = decoder_b_n113; // (signal)
  /* t48_core.vhd:209:10  */
  assign p2_read_reg_s = decoder_b_n148; // (signal)
  /* t48_core.vhd:210:10  */
  assign p2_read_exp_s = decoder_b_n149; // (signal)
  /* t48_core.vhd:211:10  */
  assign p2_output_pch_s = decoder_b_n150; // (signal)
  /* t48_core.vhd:212:10  */
  assign p2_data_s = use_p2_p2_b_n326; // (signal)
  /* t48_core.vhd:215:10  */
  assign pm_write_pcl_s = decoder_b_n114; // (signal)
  /* t48_core.vhd:216:10  */
  assign pm_read_pcl_s = decoder_b_n115; // (signal)
  /* t48_core.vhd:217:10  */
  assign pm_write_pch_s = decoder_b_n116; // (signal)
  /* t48_core.vhd:218:10  */
  assign pm_read_pch_s = decoder_b_n117; // (signal)
  /* t48_core.vhd:219:10  */
  assign pm_read_pmem_s = decoder_b_n118; // (signal)
  /* t48_core.vhd:220:10  */
  assign pm_inc_pc_s = decoder_b_n151; // (signal)
  /* t48_core.vhd:221:10  */
  assign pm_write_pmem_addr_s = decoder_b_n152; // (signal)
  /* t48_core.vhd:222:10  */
  assign pm_data_s = pmem_ctrl_b_n339; // (signal)
  /* t48_core.vhd:223:10  */
  assign pm_addr_type_s = decoder_b_n153; // (signal)
  /* t48_core.vhd:224:10  */
  assign pmem_addr_s = pmem_ctrl_b_n340; // (signal)
  /* t48_core.vhd:227:10  */
  assign psw_read_psw_s = decoder_b_n119; // (signal)
  /* t48_core.vhd:228:10  */
  assign psw_read_sp_s = decoder_b_n120; // (signal)
  /* t48_core.vhd:229:10  */
  assign psw_write_psw_s = decoder_b_n121; // (signal)
  /* t48_core.vhd:230:10  */
  assign psw_write_sp_s = decoder_b_n122; // (signal)
  /* t48_core.vhd:231:10  */
  assign psw_carry_s = psw_b_n346; // (signal)
  /* t48_core.vhd:232:10  */
  assign psw_aux_carry_s = psw_b_n347; // (signal)
  /* t48_core.vhd:233:10  */
  assign psw_f0_s = psw_b_n348; // (signal)
  /* t48_core.vhd:234:10  */
  assign psw_bs_s = psw_b_n349; // (signal)
  /* t48_core.vhd:235:10  */
  assign psw_special_data_s = decoder_b_n154; // (signal)
  /* t48_core.vhd:236:10  */
  assign psw_inc_stackp_s = decoder_b_n155; // (signal)
  /* t48_core.vhd:237:10  */
  assign psw_dec_stackp_s = decoder_b_n156; // (signal)
  /* t48_core.vhd:238:10  */
  assign psw_write_carry_s = decoder_b_n157; // (signal)
  /* t48_core.vhd:239:10  */
  assign psw_write_aux_carry_s = decoder_b_n158; // (signal)
  /* t48_core.vhd:240:10  */
  assign psw_write_f0_s = decoder_b_n159; // (signal)
  /* t48_core.vhd:241:10  */
  assign psw_write_bs_s = decoder_b_n160; // (signal)
  /* t48_core.vhd:242:10  */
  assign psw_data_s = psw_b_n345; // (signal)
  /* t48_core.vhd:245:10  */
  assign tim_overflow_s = n316_o; // (signal)
  /* t48_core.vhd:246:10  */
  assign tim_of_s = use_timer_timer_b_n304; // (signal)
  /* t48_core.vhd:247:10  */
  assign tim_read_timer_s = decoder_b_n142; // (signal)
  /* t48_core.vhd:248:10  */
  assign tim_write_timer_s = decoder_b_n143; // (signal)
  /* t48_core.vhd:249:10  */
  assign tim_start_t_s = decoder_b_n144; // (signal)
  /* t48_core.vhd:250:10  */
  assign tim_start_cnt_s = decoder_b_n145; // (signal)
  /* t48_core.vhd:251:10  */
  assign tim_stop_tcnt_s = decoder_b_n146; // (signal)
  /* t48_core.vhd:252:10  */
  assign tim_data_s = use_timer_timer_b_n303; // (signal)
  /* t48_pack-p.vhd:75:5  */
  assign n26_o = xtal_en_i ? 1'b1 : 1'b0;
  /* t48_pack-p.vhd:75:5  */
  assign n34_o = en_clk_i ? 1'b1 : 1'b0;
  /* t48_core.vhd:290:29  */
  assign alu_b_n35 = alu_b_data_o; // (signal)
  /* t48_core.vhd:296:29  */
  assign alu_b_n36 = alu_b_carry_o; // (signal)
  /* t48_core.vhd:297:29  */
  assign alu_b_n37 = alu_b_aux_carry_o; // (signal)
  /* t48_core.vhd:301:29  */
  assign alu_b_n38 = alu_b_da_overflow_o; // (signal)
  /* t48_core.vhd:284:3  */
  t48_alu alu_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_accu_i(alu_write_accu_s),
    .write_shadow_i(alu_write_shadow_s),
    .write_temp_reg_i(alu_write_temp_reg_s),
    .read_alu_i(alu_read_alu_s),
    .carry_i(psw_carry_s),
    .alu_op_i(alu_op_s),
    .use_carry_i(alu_use_carry_s),
    .da_high_i(alu_da_high_s),
    .accu_low_i(alu_accu_low_s),
    .p06_temp_reg_i(alu_p06_temp_reg_s),
    .p60_temp_reg_i(alu_p60_temp_reg_s),
    .data_o(alu_b_data_o),
    .carry_o(alu_b_carry_o),
    .aux_carry_o(alu_b_aux_carry_o),
    .da_overflow_o(alu_b_da_overflow_o));
  /* t48_core.vhd:318:21  */
  assign bus_mux_b_n47 = bus_mux_b_data_o; // (signal)
  /* t48_core.vhd:307:3  */
  t48_bus_mux bus_mux_b (
    .alu_data_i(alu_data_s),
    .bus_data_i(bus_data_s),
    .dec_data_i(dec_data_s),
    .dm_data_i(dm_data_s),
    .pm_data_i(pm_data_s),
    .p1_data_i(p1_data_s),
    .p2_data_i(p2_data_s),
    .psw_data_i(psw_data_s),
    .tim_data_i(tim_data_s),
    .data_o(bus_mux_b_data_o));
  /* t48_core.vhd:331:25  */
  assign clock_ctrl_b_n50 = clock_ctrl_b_xtal3_o; // (signal)
  /* t48_core.vhd:332:25  */
  assign clock_ctrl_b_n51 = clock_ctrl_b_t0_o; // (signal)
  /* t48_core.vhd:338:25  */
  assign clock_ctrl_b_n52 = clock_ctrl_b_mstate_o; // (signal)
  /* t48_core.vhd:339:25  */
  assign clock_ctrl_b_n53 = clock_ctrl_b_second_cycle_o; // (signal)
  /* t48_core.vhd:340:25  */
  assign clock_ctrl_b_n54 = clock_ctrl_b_ale_o; // (signal)
  /* t48_core.vhd:341:25  */
  assign clock_ctrl_b_n55 = clock_ctrl_b_psen_o; // (signal)
  /* t48_core.vhd:342:25  */
  assign clock_ctrl_b_n56 = clock_ctrl_b_prog_o; // (signal)
  /* t48_core.vhd:343:25  */
  assign clock_ctrl_b_n57 = clock_ctrl_b_rd_o; // (signal)
  /* t48_core.vhd:344:25  */
  assign clock_ctrl_b_n58 = clock_ctrl_b_wr_o; // (signal)
  /* t48_core.vhd:321:3  */
  t48_clock_ctrl_1 clock_ctrl_b (
    .clk_i(clk_i),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_s),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .multi_cycle_i(clk_multi_cycle_s),
    .assert_psen_i(clk_assert_psen_s),
    .assert_prog_i(clk_assert_prog_s),
    .assert_rd_i(clk_assert_rd_s),
    .assert_wr_i(clk_assert_wr_s),
    .xtal3_o(clock_ctrl_b_xtal3_o),
    .t0_o(clock_ctrl_b_t0_o),
    .mstate_o(clock_ctrl_b_mstate_o),
    .second_cycle_o(clock_ctrl_b_second_cycle_o),
    .ale_o(clock_ctrl_b_ale_o),
    .psen_o(clock_ctrl_b_psen_o),
    .prog_o(clock_ctrl_b_prog_o),
    .rd_o(clock_ctrl_b_rd_o),
    .wr_o(clock_ctrl_b_wr_o));
  /* t48_core.vhd:354:25  */
  assign cond_branch_b_n77 = cond_branch_b_take_branch_o; // (signal)
  /* t48_core.vhd:347:3  */
  t48_cond_branch cond_branch_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .compute_take_i(cnd_compute_take_s),
    .branch_cond_i(cnd_branch_cond_s),
    .accu_i(alu_data_s),
    .t0_i(t0_s),
    .t1_i(t1_s),
    .int_n_i(int_n_i),
    .f0_i(psw_f0_s),
    .f1_i(cnd_f1_s),
    .tf_i(cnd_tf_s),
    .carry_i(psw_carry_s),
    .ibf_i(n78_o),
    .obf_i(n79_o),
    .comp_value_i(cnd_comp_value_s),
    .take_branch_o(cond_branch_b_take_branch_o));
  /* t48_core.vhd:374:25  */
  assign use_db_bus_db_bus_b_n82 = use_db_bus_db_bus_b_data_o; // (signal)
  /* t48_core.vhd:379:36  */
  assign n83_o = pmem_addr_s[7:0];
  /* t48_core.vhd:381:25  */
  assign use_db_bus_db_bus_b_n84 = use_db_bus_db_bus_b_db_o; // (signal)
  /* t48_core.vhd:382:25  */
  assign use_db_bus_db_bus_b_n85 = use_db_bus_db_bus_b_db_dir_o; // (signal)
  /* t48_core.vhd:367:5  */
  t48_db_bus use_db_bus_db_bus_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .ea_i(ea_i),
    .data_i(t48_data_s),
    .write_bus_i(bus_write_bus_s),
    .read_bus_i(bus_read_bus_s),
    .output_pcl_i(bus_output_pcl_s),
    .bidir_bus_i(bus_bidir_bus_s),
    .pcl_i(n83_o),
    .db_i(db_i),
    .data_o(use_db_bus_db_bus_b_data_o),
    .db_o(use_db_bus_db_bus_b_db_o),
    .db_dir_o(use_db_bus_db_bus_b_db_dir_o));
  /* t48_core.vhd:405:33  */
  assign decoder_b_n92 = decoder_b_t0_dir_o; // (signal)
  /* t48_core.vhd:407:33  */
  assign decoder_b_n93 = decoder_b_data_o; // (signal)
  /* t48_core.vhd:408:33  */
  assign decoder_b_n94 = decoder_b_alu_write_accu_o; // (signal)
  /* t48_core.vhd:409:33  */
  assign decoder_b_n95 = decoder_b_alu_write_shadow_o; // (signal)
  /* t48_core.vhd:410:33  */
  assign decoder_b_n96 = decoder_b_alu_write_temp_reg_o; // (signal)
  /* t48_core.vhd:411:33  */
  assign decoder_b_n97 = decoder_b_alu_read_alu_o; // (signal)
  /* t48_core.vhd:412:33  */
  assign decoder_b_n98 = decoder_b_bus_write_bus_o; // (signal)
  /* t48_core.vhd:413:33  */
  assign decoder_b_n99 = decoder_b_bus_read_bus_o; // (signal)
  /* t48_core.vhd:414:33  */
  assign decoder_b_n106 = decoder_b_dm_write_dmem_addr_o; // (signal)
  /* t48_core.vhd:415:33  */
  assign decoder_b_n107 = decoder_b_dm_write_dmem_o; // (signal)
  /* t48_core.vhd:416:33  */
  assign decoder_b_n108 = decoder_b_dm_read_dmem_o; // (signal)
  /* t48_core.vhd:417:33  */
  assign decoder_b_n109 = decoder_b_p1_write_p1_o; // (signal)
  /* t48_core.vhd:418:33  */
  assign decoder_b_n110 = decoder_b_p1_read_p1_o; // (signal)
  /* t48_core.vhd:420:33  */
  assign decoder_b_n111 = decoder_b_p2_write_p2_o; // (signal)
  /* t48_core.vhd:421:33  */
  assign decoder_b_n112 = decoder_b_p2_write_exp_o; // (signal)
  /* t48_core.vhd:422:33  */
  assign decoder_b_n113 = decoder_b_p2_read_p2_o; // (signal)
  /* t48_core.vhd:419:33  */
  assign decoder_b_n114 = decoder_b_pm_write_pcl_o; // (signal)
  /* t48_core.vhd:423:33  */
  assign decoder_b_n115 = decoder_b_pm_read_pcl_o; // (signal)
  /* t48_core.vhd:424:33  */
  assign decoder_b_n116 = decoder_b_pm_write_pch_o; // (signal)
  /* t48_core.vhd:425:33  */
  assign decoder_b_n117 = decoder_b_pm_read_pch_o; // (signal)
  /* t48_core.vhd:426:33  */
  assign decoder_b_n118 = decoder_b_pm_read_pmem_o; // (signal)
  /* t48_core.vhd:427:33  */
  assign decoder_b_n119 = decoder_b_psw_read_psw_o; // (signal)
  /* t48_core.vhd:428:33  */
  assign decoder_b_n120 = decoder_b_psw_read_sp_o; // (signal)
  /* t48_core.vhd:429:33  */
  assign decoder_b_n121 = decoder_b_psw_write_psw_o; // (signal)
  /* t48_core.vhd:430:33  */
  assign decoder_b_n122 = decoder_b_psw_write_sp_o; // (signal)
  /* t48_core.vhd:432:33  */
  assign decoder_b_n123 = decoder_b_alu_op_o; // (signal)
  /* t48_core.vhd:434:33  */
  assign decoder_b_n124 = decoder_b_alu_da_high_o; // (signal)
  /* t48_core.vhd:436:33  */
  assign decoder_b_n125 = decoder_b_alu_accu_low_o; // (signal)
  /* t48_core.vhd:437:33  */
  assign decoder_b_n126 = decoder_b_alu_p06_temp_reg_o; // (signal)
  /* t48_core.vhd:438:33  */
  assign decoder_b_n127 = decoder_b_alu_p60_temp_reg_o; // (signal)
  /* t48_core.vhd:433:33  */
  assign decoder_b_n128 = decoder_b_alu_use_carry_o; // (signal)
  /* t48_core.vhd:439:33  */
  assign decoder_b_n129 = decoder_b_bus_output_pcl_o; // (signal)
  /* t48_core.vhd:440:33  */
  assign decoder_b_n130 = decoder_b_bus_bidir_bus_o; // (signal)
  /* t48_core.vhd:441:33  */
  assign decoder_b_n131 = decoder_b_clk_multi_cycle_o; // (signal)
  /* t48_core.vhd:442:33  */
  assign decoder_b_n132 = decoder_b_clk_assert_psen_o; // (signal)
  /* t48_core.vhd:443:33  */
  assign decoder_b_n133 = decoder_b_clk_assert_prog_o; // (signal)
  /* t48_core.vhd:444:33  */
  assign decoder_b_n134 = decoder_b_clk_assert_rd_o; // (signal)
  /* t48_core.vhd:445:33  */
  assign decoder_b_n135 = decoder_b_clk_assert_wr_o; // (signal)
  /* t48_core.vhd:448:33  */
  assign decoder_b_n136 = decoder_b_cnd_compute_take_o; // (signal)
  /* t48_core.vhd:449:33  */
  assign decoder_b_n137 = decoder_b_cnd_branch_cond_o; // (signal)
  /* t48_core.vhd:451:33  */
  assign decoder_b_n138 = decoder_b_cnd_comp_value_o; // (signal)
  /* t48_core.vhd:452:33  */
  assign decoder_b_n139 = decoder_b_cnd_f1_o; // (signal)
  /* t48_core.vhd:453:33  */
  assign decoder_b_n140 = decoder_b_cnd_tf_o; // (signal)
  /* t48_core.vhd:454:33  */
  assign decoder_b_n141 = decoder_b_dm_addr_type_o; // (signal)
  /* t48_core.vhd:455:33  */
  assign decoder_b_n142 = decoder_b_tim_read_timer_o; // (signal)
  /* t48_core.vhd:456:33  */
  assign decoder_b_n143 = decoder_b_tim_write_timer_o; // (signal)
  /* t48_core.vhd:457:33  */
  assign decoder_b_n144 = decoder_b_tim_start_t_o; // (signal)
  /* t48_core.vhd:458:33  */
  assign decoder_b_n145 = decoder_b_tim_start_cnt_o; // (signal)
  /* t48_core.vhd:459:33  */
  assign decoder_b_n146 = decoder_b_tim_stop_tcnt_o; // (signal)
  /* t48_core.vhd:460:33  */
  assign decoder_b_n147 = decoder_b_p1_read_reg_o; // (signal)
  /* t48_core.vhd:461:33  */
  assign decoder_b_n148 = decoder_b_p2_read_reg_o; // (signal)
  /* t48_core.vhd:462:33  */
  assign decoder_b_n149 = decoder_b_p2_read_exp_o; // (signal)
  /* t48_core.vhd:463:33  */
  assign decoder_b_n150 = decoder_b_p2_output_pch_o; // (signal)
  /* t48_core.vhd:464:33  */
  assign decoder_b_n151 = decoder_b_pm_inc_pc_o; // (signal)
  /* t48_core.vhd:465:33  */
  assign decoder_b_n152 = decoder_b_pm_write_pmem_addr_o; // (signal)
  /* t48_core.vhd:466:33  */
  assign decoder_b_n153 = decoder_b_pm_addr_type_o; // (signal)
  /* t48_core.vhd:467:33  */
  assign decoder_b_n154 = decoder_b_psw_special_data_o; // (signal)
  /* t48_core.vhd:471:33  */
  assign decoder_b_n155 = decoder_b_psw_inc_stackp_o; // (signal)
  /* t48_core.vhd:472:33  */
  assign decoder_b_n156 = decoder_b_psw_dec_stackp_o; // (signal)
  /* t48_core.vhd:473:33  */
  assign decoder_b_n157 = decoder_b_psw_write_carry_o; // (signal)
  /* t48_core.vhd:474:33  */
  assign decoder_b_n158 = decoder_b_psw_write_aux_carry_o; // (signal)
  /* t48_core.vhd:475:33  */
  assign decoder_b_n159 = decoder_b_psw_write_f0_o; // (signal)
  /* t48_core.vhd:476:33  */
  assign decoder_b_n160 = decoder_b_psw_write_bs_o; // (signal)
  /* t48_core.vhd:392:3  */
  t48_decoder_1_0_0 decoder_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_s),
    .ea_i(ea_i),
    .ale_i(ale_s),
    .int_n_i(int_n_i),
    .data_i(t48_data_s),
    .bus_set_f1_i(n100_o),
    .bus_clear_f1_i(n101_o),
    .alu_carry_i(alu_carry_s),
    .alu_da_overflow_i(alu_da_overflow_s),
    .clk_mstate_i(clk_mstate_s),
    .clk_second_cycle_i(clk_second_cycle_s),
    .cnd_take_branch_i(cnd_take_branch_s),
    .psw_carry_i(psw_carry_s),
    .psw_aux_carry_i(psw_aux_carry_s),
    .psw_f0_i(psw_f0_s),
    .tim_overflow_i(tim_overflow_s),
    .t0_dir_o(decoder_b_t0_dir_o),
    .data_o(decoder_b_data_o),
    .alu_write_accu_o(decoder_b_alu_write_accu_o),
    .alu_write_shadow_o(decoder_b_alu_write_shadow_o),
    .alu_write_temp_reg_o(decoder_b_alu_write_temp_reg_o),
    .alu_read_alu_o(decoder_b_alu_read_alu_o),
    .bus_write_bus_o(decoder_b_bus_write_bus_o),
    .bus_read_bus_o(decoder_b_bus_read_bus_o),
    .bus_ibf_int_o(),
    .bus_en_dma_o(),
    .bus_en_flags_o(),
    .bus_write_sts_o(),
    .dm_write_dmem_addr_o(decoder_b_dm_write_dmem_addr_o),
    .dm_write_dmem_o(decoder_b_dm_write_dmem_o),
    .dm_read_dmem_o(decoder_b_dm_read_dmem_o),
    .p1_write_p1_o(decoder_b_p1_write_p1_o),
    .p1_read_p1_o(decoder_b_p1_read_p1_o),
    .p2_write_p2_o(decoder_b_p2_write_p2_o),
    .p2_write_exp_o(decoder_b_p2_write_exp_o),
    .p2_read_p2_o(decoder_b_p2_read_p2_o),
    .p2_read_exp_o(decoder_b_p2_read_exp_o),
    .pm_write_pcl_o(decoder_b_pm_write_pcl_o),
    .pm_read_pcl_o(decoder_b_pm_read_pcl_o),
    .pm_write_pch_o(decoder_b_pm_write_pch_o),
    .pm_read_pch_o(decoder_b_pm_read_pch_o),
    .pm_read_pmem_o(decoder_b_pm_read_pmem_o),
    .psw_read_psw_o(decoder_b_psw_read_psw_o),
    .psw_read_sp_o(decoder_b_psw_read_sp_o),
    .psw_write_psw_o(decoder_b_psw_write_psw_o),
    .psw_write_sp_o(decoder_b_psw_write_sp_o),
    .alu_op_o(decoder_b_alu_op_o),
    .alu_use_carry_o(decoder_b_alu_use_carry_o),
    .alu_da_high_o(decoder_b_alu_da_high_o),
    .alu_accu_low_o(decoder_b_alu_accu_low_o),
    .alu_p06_temp_reg_o(decoder_b_alu_p06_temp_reg_o),
    .alu_p60_temp_reg_o(decoder_b_alu_p60_temp_reg_o),
    .bus_output_pcl_o(decoder_b_bus_output_pcl_o),
    .bus_bidir_bus_o(decoder_b_bus_bidir_bus_o),
    .clk_multi_cycle_o(decoder_b_clk_multi_cycle_o),
    .clk_assert_psen_o(decoder_b_clk_assert_psen_o),
    .clk_assert_prog_o(decoder_b_clk_assert_prog_o),
    .clk_assert_rd_o(decoder_b_clk_assert_rd_o),
    .clk_assert_wr_o(decoder_b_clk_assert_wr_o),
    .cnd_compute_take_o(decoder_b_cnd_compute_take_o),
    .cnd_branch_cond_o(decoder_b_cnd_branch_cond_o),
    .cnd_comp_value_o(decoder_b_cnd_comp_value_o),
    .cnd_f1_o(decoder_b_cnd_f1_o),
    .cnd_tf_o(decoder_b_cnd_tf_o),
    .dm_addr_type_o(decoder_b_dm_addr_type_o),
    .p1_read_reg_o(decoder_b_p1_read_reg_o),
    .p2_read_reg_o(decoder_b_p2_read_reg_o),
    .p2_output_pch_o(decoder_b_p2_output_pch_o),
    .pm_inc_pc_o(decoder_b_pm_inc_pc_o),
    .pm_write_pmem_addr_o(decoder_b_pm_write_pmem_addr_o),
    .pm_addr_type_o(decoder_b_pm_addr_type_o),
    .psw_special_data_o(decoder_b_psw_special_data_o),
    .psw_inc_stackp_o(decoder_b_psw_inc_stackp_o),
    .psw_dec_stackp_o(decoder_b_psw_dec_stackp_o),
    .psw_write_carry_o(decoder_b_psw_write_carry_o),
    .psw_write_aux_carry_o(decoder_b_psw_write_aux_carry_o),
    .psw_write_f0_o(decoder_b_psw_write_f0_o),
    .psw_write_bs_o(decoder_b_psw_write_bs_o),
    .tim_read_timer_o(decoder_b_tim_read_timer_o),
    .tim_write_timer_o(decoder_b_tim_write_timer_o),
    .tim_start_t_o(decoder_b_tim_start_t_o),
    .tim_start_cnt_o(decoder_b_tim_start_cnt_o),
    .tim_stop_tcnt_o(decoder_b_tim_stop_tcnt_o));
  /* t48_core.vhd:491:28  */
  assign dmem_ctrl_b_n291 = dmem_ctrl_b_data_o; // (signal)
  /* t48_core.vhd:493:28  */
  assign dmem_ctrl_b_n292 = dmem_ctrl_b_dmem_addr_o; // (signal)
  /* t48_core.vhd:494:28  */
  assign dmem_ctrl_b_n293 = dmem_ctrl_b_dmem_we_o; // (signal)
  /* t48_core.vhd:495:28  */
  assign dmem_ctrl_b_n294 = dmem_ctrl_b_dmem_data_o; // (signal)
  /* t48_core.vhd:480:3  */
  t48_dmem_ctrl dmem_ctrl_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_dmem_addr_i(dm_write_dmem_addr_s),
    .write_dmem_i(dm_write_dmem_s),
    .read_dmem_i(dm_read_dmem_s),
    .addr_type_i(dm_addr_type_s),
    .bank_select_i(psw_bs_s),
    .dmem_data_i(dmem_data_i),
    .data_o(dmem_ctrl_b_data_o),
    .dmem_addr_o(dmem_ctrl_b_dmem_addr_o),
    .dmem_we_o(dmem_ctrl_b_dmem_we_o),
    .dmem_data_o(dmem_ctrl_b_dmem_data_o));
  /* t48_core.vhd:510:26  */
  assign use_timer_timer_b_n303 = use_timer_timer_b_data_o; // (signal)
  /* t48_core.vhd:516:26  */
  assign use_timer_timer_b_n304 = use_timer_timer_b_overflow_o; // (signal)
  /* t48_core.vhd:499:5  */
  t48_timer_4 use_timer_timer_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .t1_i(t1_s),
    .clk_mstate_i(clk_mstate_s),
    .data_i(t48_data_s),
    .read_timer_i(tim_read_timer_s),
    .write_timer_i(tim_write_timer_s),
    .start_t_i(tim_start_t_s),
    .start_cnt_i(tim_start_cnt_s),
    .stop_tcnt_i(tim_stop_tcnt_s),
    .data_o(use_timer_timer_b_data_o),
    .overflow_o(use_timer_timer_b_overflow_o));
  /* t48_pack-p.vhd:75:5  */
  assign n316_o = tim_of_s ? 1'b1 : 1'b0;
  /* t48_core.vhd:534:25  */
  assign use_p1_p1_b_n317 = use_p1_p1_b_data_o; // (signal)
  /* t48_core.vhd:539:25  */
  assign use_p1_p1_b_n318 = use_p1_p1_b_p1_o; // (signal)
  /* t48_core.vhd:540:25  */
  assign use_p1_p1_b_n319 = use_p1_p1_b_p1_low_imp_o; // (signal)
  /* t48_core.vhd:528:5  */
  t48_p1 use_p1_p1_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_p1_i(p1_write_p1_s),
    .read_p1_i(p1_read_p1_s),
    .read_reg_i(p1_read_reg_s),
    .p1_i(p1_i),
    .data_o(use_p1_p1_b_data_o),
    .p1_o(use_p1_p1_b_p1_o),
    .p1_low_imp_o(use_p1_p1_b_p1_low_imp_o));
  /* t48_core.vhd:559:26  */
  assign use_p2_p2_b_n326 = use_p2_p2_b_data_o; // (signal)
  /* t48_core.vhd:566:37  */
  assign n327_o = pmem_addr_s[11:8];
  /* t48_core.vhd:568:26  */
  assign use_p2_p2_b_n328 = use_p2_p2_b_p2_o; // (signal)
  /* t48_core.vhd:569:26  */
  assign use_p2_p2_b_n329 = use_p2_p2_b_p2l_low_imp_o; // (signal)
  /* t48_core.vhd:570:26  */
  assign use_p2_p2_b_n330 = use_p2_p2_b_p2h_low_imp_o; // (signal)
  /* t48_core.vhd:551:5  */
  t48_p2 use_p2_p2_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .xtal_i(xtal_i),
    .xtal_en_i(xtal_en_s),
    .data_i(t48_data_s),
    .write_p2_i(p2_write_p2_s),
    .write_exp_i(p2_write_exp_s),
    .read_p2_i(p2_read_p2_s),
    .read_reg_i(p2_read_reg_s),
    .read_exp_i(p2_read_exp_s),
    .output_pch_i(p2_output_pch_s),
    .pch_i(n327_o),
    .p2_i(p2_i),
    .data_o(use_p2_p2_b_data_o),
    .p2_o(use_p2_p2_b_p2_o),
    .p2l_low_imp_o(use_p2_p2_b_p2l_low_imp_o),
    .p2h_low_imp_o(use_p2_p2_b_p2h_low_imp_o));
  /* t48_core.vhd:587:28  */
  assign pmem_ctrl_b_n339 = pmem_ctrl_b_data_o; // (signal)
  /* t48_core.vhd:596:28  */
  assign pmem_ctrl_b_n340 = pmem_ctrl_b_pmem_addr_o; // (signal)
  /* t48_core.vhd:581:3  */
  t48_pmem_ctrl pmem_ctrl_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .write_pcl_i(pm_write_pcl_s),
    .read_pcl_i(pm_read_pcl_s),
    .write_pch_i(pm_write_pch_s),
    .read_pch_i(pm_read_pch_s),
    .inc_pc_i(pm_inc_pc_s),
    .write_pmem_addr_i(pm_write_pmem_addr_s),
    .addr_type_i(pm_addr_type_s),
    .read_pmem_i(pm_read_pmem_s),
    .pmem_data_i(pmem_data_i),
    .data_o(pmem_ctrl_b_data_o),
    .pmem_addr_o(pmem_ctrl_b_pmem_addr_o));
  /* t48_core.vhd:606:29  */
  assign psw_b_n345 = psw_b_data_o; // (signal)
  /* t48_core.vhd:618:29  */
  assign psw_b_n346 = psw_b_carry_o; // (signal)
  /* t48_core.vhd:620:29  */
  assign psw_b_n347 = psw_b_aux_carry_o; // (signal)
  /* t48_core.vhd:621:29  */
  assign psw_b_n348 = psw_b_f0_o; // (signal)
  /* t48_core.vhd:622:29  */
  assign psw_b_n349 = psw_b_bs_o; // (signal)
  /* t48_core.vhd:600:3  */
  t48_psw psw_b (
    .clk_i(clk_i),
    .res_i(reset_i),
    .en_clk_i(en_clk_s),
    .data_i(t48_data_s),
    .read_psw_i(psw_read_psw_s),
    .read_sp_i(psw_read_sp_s),
    .write_psw_i(psw_write_psw_s),
    .write_sp_i(psw_write_sp_s),
    .special_data_i(psw_special_data_s),
    .inc_stackp_i(psw_inc_stackp_s),
    .dec_stackp_i(psw_dec_stackp_s),
    .write_carry_i(psw_write_carry_s),
    .write_aux_carry_i(psw_write_aux_carry_s),
    .write_f0_i(psw_write_f0_s),
    .write_bs_i(psw_write_bs_s),
    .aux_carry_i(alu_aux_carry_s),
    .data_o(psw_b_data_o),
    .carry_o(psw_b_carry_o),
    .aux_carry_o(psw_b_aux_carry_o),
    .f0_o(psw_b_f0_o),
    .bs_o(psw_b_bs_o));
  /* t48_pack-p.vhd:66:5  */
  assign n367_o = ale_s ? 1'b1 : 1'b0;
  /* t48_core.vhd:630:30  */
  assign n369_o = ~psen_s;
  /* t48_pack-p.vhd:66:5  */
  assign n376_o = n369_o ? 1'b1 : 1'b0;
  /* t48_core.vhd:631:30  */
  assign n378_o = ~prog_s;
  /* t48_pack-p.vhd:66:5  */
  assign n385_o = n378_o ? 1'b1 : 1'b0;
  /* t48_core.vhd:632:30  */
  assign n387_o = ~rd_s;
  /* t48_pack-p.vhd:66:5  */
  assign n394_o = n387_o ? 1'b1 : 1'b0;
  /* t48_core.vhd:633:30  */
  assign n396_o = ~wr_s;
  /* t48_pack-p.vhd:66:5  */
  assign n403_o = n396_o ? 1'b1 : 1'b0;
  /* t48_pack-p.vhd:66:5  */
  assign n411_o = xtal3_s ? 1'b1 : 1'b0;
endmodule

