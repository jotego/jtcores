module jt_gng;

	jt7641 sh5_2k(
		.d	( 4'd0 ),
		
	);
endmodule

