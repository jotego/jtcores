/*  This file is part of JTCORES.
    JTCORES program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTCORES program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTCORES.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 15-11-2025 */

module jtcal50_video(
    input               rst,
    input               clk,
    input               clk_cpu,
    input               pxl2_cen,
    input               pxl_cen,

    output              LHBL,
    output              LVBL,
    output              HS,
    output              VS,
    output              flip,
    // Palette
    output     [ 9:1]   pal_addr,
    input      [15:0]   pal_data,
    // CPU      interface
    input               cpu_rnw,
    input      [12:0]   cpu_addr,
    input      [15:0]   cpu_dout,
    input      [ 1:0]   cpu_dsn,
    input               vram_cs,
    input               vctrl_cs,
    input               vflag_cs,
    output     [15:0]   vram_dout,
    // SDRAM interface
    output     [20:2]   scr_addr,
    input      [31:0]   scr_data,
    input               scr_ok,
    output              scr_cs,

    output     [20:2]   obj_addr,
    input      [31:0]   obj_data,
    input               obj_ok,
    output              obj_cs,
    // Colours
    output     [ 4:0]   red,
    output     [ 4:0]   green,
    output     [ 4:0]   blue,
    // Test
    input      [ 3:0]   gfx_en,
    input      [ 7:0]   debug_bus,
    output     [ 7:0]   st_dout
);

wire [ 8:0] vrender, vrender1, hdump, vdump;
wire [ 8:0] scr_pxl, obj_pxl;

// Measured on PCB
// 64us per line, 8us blanking
// 17.45ms per frame, 2.05ms blanking, 512.5us sync (centered)
jtframe_vtimer #(
    .HB_END  ( 9'd0   ),
    .HB_START( 9'd384 ),
    .HS_START( 9'd416 ),
    .HS_END  ( 9'd480 ),
    .HCNT_END( 9'd511 ),
    .V_START ( 9'd000 ),
    .VS_START( 9'd252 ),
    .VS_END  ( 9'd260 ),
    .VB_START( 9'd239 ),
    .VB_END  ( 9'd271 ),
    .VCNT_END( 9'd271 )
) u_timer(
    .clk        ( clk        ),
    .pxl_cen    ( pxl_cen    ),
    .vdump      ( vdump      ),
    .vrender    ( vrender    ),
    .vrender1   ( vrender1   ),
    .H          ( hdump      ),
    .Hinit      (            ),
    .Vinit      (            ),
    .LHBL       ( LHBL       ),
    .LVBL       ( LVBL       ),
    .HS         ( HS         ),
    .VS         ( VS         )
);

jtkiwi_gfx #(.CPUW(16)) u_gfx(
    .rst        ( rst            ),
    .clk        ( clk            ),
    .clk_cpu    ( clk_cpu        ),
    .pxl_cen    ( pxl_cen        ),
    .pxl2_cen   ( pxl2_cen       ),
    // Screen
    .flip       ( flip           ),
    .LHBL       ( LHBL           ),
    .LVBL       ( LVBL           ),
    .vs         ( VS             ),
    .hs         ( HS             ),
    .vdump      ( vdump          ),
    .vrender    ( vrender        ),
    .hdump      ( hdump          ),
    // CPU interface
    .vram_cs    ( vram_cs        ),
    .vctrl_cs   ( vctrl_cs       ),
    .vflag_cs   ( vflag_cs       ),
    .cpu_addr   ( cpu_addr       ),
    .cpu_rnw    ( cpu_rnw        ),
    .cpu_dout   ( cpu_dout       ),
    .cpu_din    ( vram_dout      ),
    // 16-bit interface
    .cpu_dsn    ( cpu_dsn        ),
    // SDRAM
    .scr_addr   ( scr_addr       ),
    .scr_data   ( scr_data       ),
    .scr_ok     ( scr_ok         ),
    .scr_cs     ( scr_cs         ),

    .obj_addr   ( obj_addr       ),
    .obj_data   ( obj_data       ),
    .obj_ok     ( obj_ok         ),
    .obj_cs     ( obj_cs         ),
    // Color address to palette
    .scr_pxl    ( scr_pxl        ),
    .obj_pxl    ( obj_pxl        ),
    .debug_bus  ( debug_bus      ),
    .st_dout    ( st_dout        )
);

jtcal50_colmix u_colmix(
    .clk        ( clk            ),
    .clk_cpu    ( clk_cpu        ),
    .pxl_cen    ( pxl_cen        ),
    // Screen
    .LHBL       ( LHBL           ),
    .LVBL       ( LVBL           ),
    // RAM
    .pal_addr   ( pal_addr       ),
    .pal_data   ( pal_data       ),
    // Colour output
    .scr_pxl    ( scr_pxl        ),
    .obj_pxl    ( obj_pxl        ),
    .red        ( red            ),
    .green      ( green          ),
    .blue       ( blue           ),
    .gfx_en     ( gfx_en         ),
    .debug_bus  ( debug_bus      )
);

endmodule
