module test;

localparam W=7; //8
localparam [7:0] OFFSET='h40;

reg clk, rst;
reg [7:0] dout;
reg play;
wire signed [W-1:0] snd;

/*
initial begin
    $dumpfile("test.lxt");
    $dumpvars;
    $dumpon;
    #10000000 $finish;
end
*/

initial begin
    clk=0;
    forever #10 clk=~clk;
end

integer gain=0,exp;

initial begin
    rst  = 1;
    play = 0;
    dout=0;
    repeat (20) @(posedge clk);
    rst  = 0;
    @(posedge clk)
    play = 1;
    for(gain=0;gain<256;gain=gain+1) begin
        dout=gain[7:0];
        repeat (2) @(posedge clk);
        exp = dout[6:0] - OFFSET;
        @(posedge clk);
        if(snd!=$signed(exp[W-1:0])) begin
            $display("Bad value at rom_dout %d",dout);
            $display("output vs expected: %d <> %d",snd,exp);
            $display("FAIL");
            $finish;
        end
        if( exp[30:W-1]!={32-W{exp[31]}}) begin
            $display("Bad sign at rom_dout %d/%d",dout);
            $display("output vs expected: %d <> %d",snd,exp);
            $display("FAIL");
            $finish;
        end
    end
    $display("PASS");
    $finish;
end


jt007232_channel uut(
    .rst        ( rst     ),
    .clk        ( clk     ),
    .cen_q      ( 1'b1    ),
    .rom_start  ( 17'h0   ),
    .pre0       ( 12'hFFF ),
    .pre_sel    ( 2'b0    ),
    .loop       ( 1'b1    ),
    .play       ( play    ),
    .load       ( 1'b1    ),
    .rom_addr   (         ),
    .rom_cs     (         ),
    .rom_ok     ( 1'b1    ),
    .rom_dout   ( dout    ),
    .snd        ( snd     )
);

endmodule