localparam [8:0]
    V_START  = 9'h0F8,
    VB_START = 9'h0F8,
    VB_END   = 9'h120,
    VS_START = 9'h108,
    VS_END   = 9'h110,
    VCNT_END = 9'h1FF,
    HS_START = 9'h17f,
    HS_END   = 9'h01f,
    HB_START = 9'h160, // 288 visible, 384 total (96 pxl=HB)
    HB_END   = 9'h040;
