localparam [8:0]
    V_START  = 9'h0F8,
    VB_START = 9'h0F8,
    VB_END   = 9'h120,
    VS_START = 9'h108,
    VS_END   = 9'h110,
    VCNT_END = 9'h1FF;
