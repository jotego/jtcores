library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ccfac287",
    12 => x"86c0c54e",
    13 => x"49ccfac2",
    14 => x"48c0e7c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e7e0",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"711e4f26",
    53 => x"4966c44a",
    54 => x"c888c148",
    55 => x"997158a6",
    56 => x"ff87d602",
    57 => x"ffc348d4",
    58 => x"c4526878",
    59 => x"c1484966",
    60 => x"58a6c888",
    61 => x"ea059971",
    62 => x"1e4f2687",
    63 => x"d4ff1e73",
    64 => x"7bffc34b",
    65 => x"ffc34a6b",
    66 => x"c8496b7b",
    67 => x"c3b17232",
    68 => x"4a6b7bff",
    69 => x"b27131c8",
    70 => x"6b7bffc3",
    71 => x"7232c849",
    72 => x"c44871b1",
    73 => x"264d2687",
    74 => x"264b264c",
    75 => x"5b5e0e4f",
    76 => x"710e5d5c",
    77 => x"4cd4ff4a",
    78 => x"ffc34972",
    79 => x"c27c7199",
    80 => x"05bfc0e7",
    81 => x"66d087c8",
    82 => x"d430c948",
    83 => x"66d058a6",
    84 => x"c329d849",
    85 => x"7c7199ff",
    86 => x"d04966d0",
    87 => x"99ffc329",
    88 => x"66d07c71",
    89 => x"c329c849",
    90 => x"7c7199ff",
    91 => x"c34966d0",
    92 => x"7c7199ff",
    93 => x"29d04972",
    94 => x"7199ffc3",
    95 => x"c94b6c7c",
    96 => x"c34dfff0",
    97 => x"d005abff",
    98 => x"7cffc387",
    99 => x"8dc14b6c",
   100 => x"c387c602",
   101 => x"f002abff",
   102 => x"fe487387",
   103 => x"c01e87c7",
   104 => x"48d4ff49",
   105 => x"c178ffc3",
   106 => x"b7c8c381",
   107 => x"87f104a9",
   108 => x"731e4f26",
   109 => x"c487e71e",
   110 => x"c04bdff8",
   111 => x"f0ffc01e",
   112 => x"fd49f7c1",
   113 => x"86c487e7",
   114 => x"c005a8c1",
   115 => x"d4ff87ea",
   116 => x"78ffc348",
   117 => x"c0c0c0c1",
   118 => x"c01ec0c0",
   119 => x"e9c1f0e1",
   120 => x"87c9fd49",
   121 => x"987086c4",
   122 => x"ff87ca05",
   123 => x"ffc348d4",
   124 => x"cb48c178",
   125 => x"87e6fe87",
   126 => x"fe058bc1",
   127 => x"48c087fd",
   128 => x"1e87e6fc",
   129 => x"d4ff1e73",
   130 => x"78ffc348",
   131 => x"1ec04bd3",
   132 => x"c1f0ffc0",
   133 => x"d4fc49c1",
   134 => x"7086c487",
   135 => x"87ca0598",
   136 => x"c348d4ff",
   137 => x"48c178ff",
   138 => x"f1fd87cb",
   139 => x"058bc187",
   140 => x"c087dbff",
   141 => x"87f1fb48",
   142 => x"5c5b5e0e",
   143 => x"4cd4ff0e",
   144 => x"c687dbfd",
   145 => x"e1c01eea",
   146 => x"49c8c1f0",
   147 => x"c487defb",
   148 => x"02a8c186",
   149 => x"eafe87c8",
   150 => x"c148c087",
   151 => x"dafa87e2",
   152 => x"cf497087",
   153 => x"c699ffff",
   154 => x"c802a9ea",
   155 => x"87d3fe87",
   156 => x"cbc148c0",
   157 => x"7cffc387",
   158 => x"fc4bf1c0",
   159 => x"987087f4",
   160 => x"87ebc002",
   161 => x"ffc01ec0",
   162 => x"49fac1f0",
   163 => x"c487defa",
   164 => x"05987086",
   165 => x"ffc387d9",
   166 => x"c3496c7c",
   167 => x"7c7c7cff",
   168 => x"99c0c17c",
   169 => x"c187c402",
   170 => x"c087d548",
   171 => x"c287d148",
   172 => x"87c405ab",
   173 => x"87c848c0",
   174 => x"fe058bc1",
   175 => x"48c087fd",
   176 => x"1e87e4f9",
   177 => x"e7c21e73",
   178 => x"78c148c0",
   179 => x"d0ff4bc7",
   180 => x"fb78c248",
   181 => x"d0ff87c8",
   182 => x"c078c348",
   183 => x"d0e5c01e",
   184 => x"f949c0c1",
   185 => x"86c487c7",
   186 => x"c105a8c1",
   187 => x"abc24b87",
   188 => x"c087c505",
   189 => x"87f9c048",
   190 => x"ff058bc1",
   191 => x"f7fc87d0",
   192 => x"c4e7c287",
   193 => x"05987058",
   194 => x"1ec187cd",
   195 => x"c1f0ffc0",
   196 => x"d8f849d0",
   197 => x"ff86c487",
   198 => x"ffc348d4",
   199 => x"87fcc278",
   200 => x"58c8e7c2",
   201 => x"c248d0ff",
   202 => x"48d4ff78",
   203 => x"c178ffc3",
   204 => x"87f5f748",
   205 => x"5c5b5e0e",
   206 => x"4b710e5d",
   207 => x"eec54cc0",
   208 => x"ff4adfcd",
   209 => x"ffc348d4",
   210 => x"c3496878",
   211 => x"c005a9fe",
   212 => x"4d7087fd",
   213 => x"cc029b73",
   214 => x"1e66d087",
   215 => x"f1f54973",
   216 => x"d686c487",
   217 => x"48d0ff87",
   218 => x"c378d1c4",
   219 => x"66d07dff",
   220 => x"d488c148",
   221 => x"987058a6",
   222 => x"ff87f005",
   223 => x"ffc348d4",
   224 => x"9b737878",
   225 => x"ff87c505",
   226 => x"78d048d0",
   227 => x"c14c4ac1",
   228 => x"eefe058a",
   229 => x"f6487487",
   230 => x"731e87cb",
   231 => x"c04a711e",
   232 => x"48d4ff4b",
   233 => x"ff78ffc3",
   234 => x"c3c448d0",
   235 => x"48d4ff78",
   236 => x"7278ffc3",
   237 => x"f0ffc01e",
   238 => x"f549d1c1",
   239 => x"86c487ef",
   240 => x"d2059870",
   241 => x"1ec0c887",
   242 => x"fd4966cc",
   243 => x"86c487e6",
   244 => x"d0ff4b70",
   245 => x"7378c248",
   246 => x"87cdf548",
   247 => x"5c5b5e0e",
   248 => x"1ec00e5d",
   249 => x"c1f0ffc0",
   250 => x"c0f549c9",
   251 => x"c21ed287",
   252 => x"fc49c8e7",
   253 => x"86c887fe",
   254 => x"84c14cc0",
   255 => x"04acb7d2",
   256 => x"e7c287f8",
   257 => x"49bf97c8",
   258 => x"c199c0c3",
   259 => x"c005a9c0",
   260 => x"e7c287e7",
   261 => x"49bf97cf",
   262 => x"e7c231d0",
   263 => x"4abf97d0",
   264 => x"b17232c8",
   265 => x"97d1e7c2",
   266 => x"71b14abf",
   267 => x"ffffcf4c",
   268 => x"84c19cff",
   269 => x"e7c134ca",
   270 => x"d1e7c287",
   271 => x"c149bf97",
   272 => x"c299c631",
   273 => x"bf97d2e7",
   274 => x"2ab7c74a",
   275 => x"e7c2b172",
   276 => x"4abf97cd",
   277 => x"c29dcf4d",
   278 => x"bf97cee7",
   279 => x"ca9ac34a",
   280 => x"cfe7c232",
   281 => x"c24bbf97",
   282 => x"c2b27333",
   283 => x"bf97d0e7",
   284 => x"9bc0c34b",
   285 => x"732bb7c6",
   286 => x"c181c2b2",
   287 => x"70307148",
   288 => x"7548c149",
   289 => x"724d7030",
   290 => x"7184c14c",
   291 => x"b7c0c894",
   292 => x"87cc06ad",
   293 => x"2db734c1",
   294 => x"adb7c0c8",
   295 => x"87f4ff01",
   296 => x"c0f24874",
   297 => x"5b5e0e87",
   298 => x"f80e5d5c",
   299 => x"eeefc286",
   300 => x"c278c048",
   301 => x"c01ee6e7",
   302 => x"87defb49",
   303 => x"987086c4",
   304 => x"c087c505",
   305 => x"87cec948",
   306 => x"7ec14dc0",
   307 => x"bfdaf5c0",
   308 => x"dce8c249",
   309 => x"4bc8714a",
   310 => x"7087cfee",
   311 => x"87c20598",
   312 => x"f5c07ec0",
   313 => x"c249bfd6",
   314 => x"714af8e8",
   315 => x"f9ed4bc8",
   316 => x"05987087",
   317 => x"7ec087c2",
   318 => x"fdc0026e",
   319 => x"eceec287",
   320 => x"efc24dbf",
   321 => x"7ebf9fe4",
   322 => x"ead6c548",
   323 => x"87c705a8",
   324 => x"bfeceec2",
   325 => x"6e87ce4d",
   326 => x"d5e9ca48",
   327 => x"87c502a8",
   328 => x"f1c748c0",
   329 => x"e6e7c287",
   330 => x"f949751e",
   331 => x"86c487ec",
   332 => x"c5059870",
   333 => x"c748c087",
   334 => x"f5c087dc",
   335 => x"c249bfd6",
   336 => x"714af8e8",
   337 => x"e1ec4bc8",
   338 => x"05987087",
   339 => x"efc287c8",
   340 => x"78c148ee",
   341 => x"f5c087da",
   342 => x"c249bfda",
   343 => x"714adce8",
   344 => x"c5ec4bc8",
   345 => x"02987087",
   346 => x"c087c5c0",
   347 => x"87e6c648",
   348 => x"97e4efc2",
   349 => x"d5c149bf",
   350 => x"cdc005a9",
   351 => x"e5efc287",
   352 => x"c249bf97",
   353 => x"c002a9ea",
   354 => x"48c087c5",
   355 => x"c287c7c6",
   356 => x"bf97e6e7",
   357 => x"e9c3487e",
   358 => x"cec002a8",
   359 => x"c3486e87",
   360 => x"c002a8eb",
   361 => x"48c087c5",
   362 => x"c287ebc5",
   363 => x"bf97f1e7",
   364 => x"c0059949",
   365 => x"e7c287cc",
   366 => x"49bf97f2",
   367 => x"c002a9c2",
   368 => x"48c087c5",
   369 => x"c287cfc5",
   370 => x"bf97f3e7",
   371 => x"eaefc248",
   372 => x"484c7058",
   373 => x"efc288c1",
   374 => x"e7c258ee",
   375 => x"49bf97f4",
   376 => x"e7c28175",
   377 => x"4abf97f5",
   378 => x"a17232c8",
   379 => x"fbf3c27e",
   380 => x"c2786e48",
   381 => x"bf97f6e7",
   382 => x"58a6c848",
   383 => x"bfeeefc2",
   384 => x"87d4c202",
   385 => x"bfd6f5c0",
   386 => x"f8e8c249",
   387 => x"4bc8714a",
   388 => x"7087d7e9",
   389 => x"c5c00298",
   390 => x"c348c087",
   391 => x"efc287f8",
   392 => x"c24cbfe6",
   393 => x"c25ccff4",
   394 => x"bf97cbe8",
   395 => x"c231c849",
   396 => x"bf97cae8",
   397 => x"c249a14a",
   398 => x"bf97cce8",
   399 => x"7232d04a",
   400 => x"e8c249a1",
   401 => x"4abf97cd",
   402 => x"a17232d8",
   403 => x"9166c449",
   404 => x"bffbf3c2",
   405 => x"c3f4c281",
   406 => x"d3e8c259",
   407 => x"c84abf97",
   408 => x"d2e8c232",
   409 => x"a24bbf97",
   410 => x"d4e8c24a",
   411 => x"d04bbf97",
   412 => x"4aa27333",
   413 => x"97d5e8c2",
   414 => x"9bcf4bbf",
   415 => x"a27333d8",
   416 => x"c7f4c24a",
   417 => x"c3f4c25a",
   418 => x"8ac24abf",
   419 => x"f4c29274",
   420 => x"a17248c7",
   421 => x"87cac178",
   422 => x"97f8e7c2",
   423 => x"31c849bf",
   424 => x"97f7e7c2",
   425 => x"49a14abf",
   426 => x"59f6efc2",
   427 => x"bff2efc2",
   428 => x"c731c549",
   429 => x"29c981ff",
   430 => x"59cff4c2",
   431 => x"97fde7c2",
   432 => x"32c84abf",
   433 => x"97fce7c2",
   434 => x"4aa24bbf",
   435 => x"6e9266c4",
   436 => x"cbf4c282",
   437 => x"c3f4c25a",
   438 => x"c278c048",
   439 => x"7248fff3",
   440 => x"f4c278a1",
   441 => x"f4c248cf",
   442 => x"c278bfc3",
   443 => x"c248d3f4",
   444 => x"78bfc7f4",
   445 => x"bfeeefc2",
   446 => x"87c9c002",
   447 => x"30c44874",
   448 => x"c9c07e70",
   449 => x"cbf4c287",
   450 => x"30c448bf",
   451 => x"efc27e70",
   452 => x"786e48f2",
   453 => x"8ef848c1",
   454 => x"4c264d26",
   455 => x"4f264b26",
   456 => x"5c5b5e0e",
   457 => x"4a710e5d",
   458 => x"bfeeefc2",
   459 => x"7287cb02",
   460 => x"722bc74b",
   461 => x"9cffc14c",
   462 => x"4b7287c9",
   463 => x"4c722bc8",
   464 => x"c29cffc3",
   465 => x"83bffbf3",
   466 => x"bfd2f5c0",
   467 => x"87d902ab",
   468 => x"5bd6f5c0",
   469 => x"1ee6e7c2",
   470 => x"fdf04973",
   471 => x"7086c487",
   472 => x"87c50598",
   473 => x"e6c048c0",
   474 => x"eeefc287",
   475 => x"87d202bf",
   476 => x"91c44974",
   477 => x"81e6e7c2",
   478 => x"ffcf4d69",
   479 => x"9dffffff",
   480 => x"497487cb",
   481 => x"e7c291c2",
   482 => x"699f81e6",
   483 => x"fe48754d",
   484 => x"5e0e87c6",
   485 => x"0e5d5c5b",
   486 => x"c04d711e",
   487 => x"cf49c11e",
   488 => x"86c487d4",
   489 => x"029c4c70",
   490 => x"c287c0c1",
   491 => x"754af6ef",
   492 => x"87dbe249",
   493 => x"c0029870",
   494 => x"4a7487f1",
   495 => x"4bcb4975",
   496 => x"7087c1e3",
   497 => x"e2c00298",
   498 => x"741ec087",
   499 => x"87c7029c",
   500 => x"c048a6c4",
   501 => x"c487c578",
   502 => x"78c148a6",
   503 => x"ce4966c4",
   504 => x"86c487d4",
   505 => x"059c4c70",
   506 => x"7487c0ff",
   507 => x"e7fc2648",
   508 => x"5b5e0e87",
   509 => x"1e0e5d5c",
   510 => x"059b4b71",
   511 => x"48c087c5",
   512 => x"c887e5c1",
   513 => x"7dc04da3",
   514 => x"c70266d4",
   515 => x"9766d487",
   516 => x"87c505bf",
   517 => x"cfc148c0",
   518 => x"4966d487",
   519 => x"7087f3fd",
   520 => x"c1029c4c",
   521 => x"a4dc87c0",
   522 => x"da7d6949",
   523 => x"a3c449a4",
   524 => x"7a699f4a",
   525 => x"bfeeefc2",
   526 => x"d487d202",
   527 => x"699f49a4",
   528 => x"ffffc049",
   529 => x"d0487199",
   530 => x"c27e7030",
   531 => x"6e7ec087",
   532 => x"806a4849",
   533 => x"7bc07a70",
   534 => x"6a49a3cc",
   535 => x"49a3d079",
   536 => x"487479c0",
   537 => x"48c087c2",
   538 => x"87ecfa26",
   539 => x"5c5b5e0e",
   540 => x"4c710e5d",
   541 => x"cac1029c",
   542 => x"49a4c887",
   543 => x"c2c10269",
   544 => x"4a66d087",
   545 => x"d482496c",
   546 => x"66d05aa6",
   547 => x"efc2b94d",
   548 => x"ff4abfea",
   549 => x"719972ba",
   550 => x"e4c00299",
   551 => x"4ba4c487",
   552 => x"fbf9496b",
   553 => x"c27b7087",
   554 => x"49bfe6ef",
   555 => x"7c71816c",
   556 => x"efc2b975",
   557 => x"ff4abfea",
   558 => x"719972ba",
   559 => x"dcff0599",
   560 => x"f97c7587",
   561 => x"731e87d2",
   562 => x"9b4b711e",
   563 => x"c887c702",
   564 => x"056949a3",
   565 => x"48c087c5",
   566 => x"c287efc0",
   567 => x"4abffff3",
   568 => x"6949a3c4",
   569 => x"c289c249",
   570 => x"91bfe6ef",
   571 => x"c24aa271",
   572 => x"49bfeaef",
   573 => x"a271996b",
   574 => x"d6f5c04a",
   575 => x"1e66c85a",
   576 => x"d5ea4972",
   577 => x"7086c487",
   578 => x"cff84849",
   579 => x"5b5e0e87",
   580 => x"1e0e5d5c",
   581 => x"66d44b71",
   582 => x"732cc94c",
   583 => x"cfc1029b",
   584 => x"49a3c887",
   585 => x"c7c10269",
   586 => x"4da3d087",
   587 => x"c27d66d4",
   588 => x"49bfeaef",
   589 => x"4a6bb9ff",
   590 => x"ac717e99",
   591 => x"c087cd03",
   592 => x"a3cc7d7b",
   593 => x"49a3c44a",
   594 => x"87c2796a",
   595 => x"9c748c72",
   596 => x"4987dd02",
   597 => x"fc49731e",
   598 => x"86c487d2",
   599 => x"c74966d4",
   600 => x"cb0299ff",
   601 => x"e6e7c287",
   602 => x"fd49731e",
   603 => x"86c487d8",
   604 => x"87e4f626",
   605 => x"5c5b5e0e",
   606 => x"86f00e5d",
   607 => x"c059a6d0",
   608 => x"cc4b66e4",
   609 => x"87ca0266",
   610 => x"7080c848",
   611 => x"05bf6e7e",
   612 => x"48c087c5",
   613 => x"cc87ecc3",
   614 => x"84d04c66",
   615 => x"a6c44973",
   616 => x"c4786c48",
   617 => x"80c48166",
   618 => x"c878bf6e",
   619 => x"c606a966",
   620 => x"66c44987",
   621 => x"c04b7189",
   622 => x"c401abb7",
   623 => x"c2c34887",
   624 => x"4866c487",
   625 => x"7098ffc7",
   626 => x"c1026e7e",
   627 => x"c0c887c9",
   628 => x"71896e49",
   629 => x"e6e7c24a",
   630 => x"73856e4d",
   631 => x"c106aab7",
   632 => x"49724a87",
   633 => x"8066c448",
   634 => x"8b727c70",
   635 => x"718ac149",
   636 => x"87d90299",
   637 => x"4866e0c0",
   638 => x"e0c05015",
   639 => x"80c14866",
   640 => x"58a6e4c0",
   641 => x"8ac14972",
   642 => x"e7059971",
   643 => x"d01ec187",
   644 => x"d7f94966",
   645 => x"c086c487",
   646 => x"c106abb7",
   647 => x"e0c087e3",
   648 => x"ffc74d66",
   649 => x"c006abb7",
   650 => x"1e7587e2",
   651 => x"fa4966d0",
   652 => x"c0c887d4",
   653 => x"c8486c85",
   654 => x"7c7080c0",
   655 => x"c18bc0c8",
   656 => x"4966d41e",
   657 => x"c887e5f8",
   658 => x"87eec086",
   659 => x"1ee6e7c2",
   660 => x"f94966d0",
   661 => x"86c487f0",
   662 => x"4ae6e7c2",
   663 => x"6c484973",
   664 => x"737c7080",
   665 => x"718bc149",
   666 => x"87ce0299",
   667 => x"c17d9712",
   668 => x"c1497385",
   669 => x"0599718b",
   670 => x"b7c087f2",
   671 => x"e1fe01ab",
   672 => x"f048c187",
   673 => x"87d0f28e",
   674 => x"5c5b5e0e",
   675 => x"4b710e5d",
   676 => x"87c7029b",
   677 => x"6d4da3c8",
   678 => x"ff87c505",
   679 => x"87fdc048",
   680 => x"6c4ca3d0",
   681 => x"99ffc749",
   682 => x"6c87d805",
   683 => x"c187c902",
   684 => x"f649731e",
   685 => x"86c487f6",
   686 => x"1ee6e7c2",
   687 => x"c5f84973",
   688 => x"6c86c487",
   689 => x"04aa6d4a",
   690 => x"48ff87c4",
   691 => x"a2c187cf",
   692 => x"c749727c",
   693 => x"e7c299ff",
   694 => x"699781e6",
   695 => x"87f8f048",
   696 => x"711e731e",
   697 => x"c0029b4b",
   698 => x"f4c287e4",
   699 => x"4a735bd3",
   700 => x"efc28ac2",
   701 => x"9249bfe6",
   702 => x"bffff3c2",
   703 => x"c2807248",
   704 => x"7158d7f4",
   705 => x"c230c448",
   706 => x"c058f6ef",
   707 => x"f4c287ed",
   708 => x"f4c248cf",
   709 => x"c278bfc3",
   710 => x"c248d3f4",
   711 => x"78bfc7f4",
   712 => x"bfeeefc2",
   713 => x"c287c902",
   714 => x"49bfe6ef",
   715 => x"87c731c4",
   716 => x"bfcbf4c2",
   717 => x"c231c449",
   718 => x"ef59f6ef",
   719 => x"5e0e87de",
   720 => x"710e5c5b",
   721 => x"724bc04a",
   722 => x"e1c0029a",
   723 => x"49a2da87",
   724 => x"c24b699f",
   725 => x"02bfeeef",
   726 => x"a2d487cf",
   727 => x"49699f49",
   728 => x"ffffc04c",
   729 => x"c234d09c",
   730 => x"744cc087",
   731 => x"4973b349",
   732 => x"ee87edfd",
   733 => x"5e0e87e4",
   734 => x"0e5d5c5b",
   735 => x"4a7186f4",
   736 => x"9a727ec0",
   737 => x"c287d802",
   738 => x"c048e2e7",
   739 => x"dae7c278",
   740 => x"d3f4c248",
   741 => x"e7c278bf",
   742 => x"f4c248de",
   743 => x"c278bfcf",
   744 => x"c048c3f0",
   745 => x"f2efc250",
   746 => x"e7c249bf",
   747 => x"714abfe2",
   748 => x"cac403aa",
   749 => x"cf497287",
   750 => x"eac00599",
   751 => x"d2f5c087",
   752 => x"dae7c248",
   753 => x"e7c278bf",
   754 => x"e7c21ee6",
   755 => x"c249bfda",
   756 => x"c148dae7",
   757 => x"ff7178a1",
   758 => x"c487ffde",
   759 => x"cef5c086",
   760 => x"e6e7c248",
   761 => x"c087cc78",
   762 => x"48bfcef5",
   763 => x"c080e0c0",
   764 => x"c258d2f5",
   765 => x"48bfe2e7",
   766 => x"e7c280c1",
   767 => x"4e2758e6",
   768 => x"bf00000d",
   769 => x"9d4dbf97",
   770 => x"87e3c202",
   771 => x"02ade5c3",
   772 => x"c087dcc2",
   773 => x"4bbfcef5",
   774 => x"1149a3cb",
   775 => x"05accf4c",
   776 => x"7587d2c1",
   777 => x"c199df49",
   778 => x"c291cd89",
   779 => x"c181f6ef",
   780 => x"51124aa3",
   781 => x"124aa3c3",
   782 => x"4aa3c551",
   783 => x"a3c75112",
   784 => x"c951124a",
   785 => x"51124aa3",
   786 => x"124aa3ce",
   787 => x"4aa3d051",
   788 => x"a3d25112",
   789 => x"d451124a",
   790 => x"51124aa3",
   791 => x"124aa3d6",
   792 => x"4aa3d851",
   793 => x"a3dc5112",
   794 => x"de51124a",
   795 => x"51124aa3",
   796 => x"fac07ec1",
   797 => x"c8497487",
   798 => x"ebc00599",
   799 => x"d0497487",
   800 => x"87d10599",
   801 => x"c00266dc",
   802 => x"497387cb",
   803 => x"700f66dc",
   804 => x"d3c00298",
   805 => x"c0056e87",
   806 => x"efc287c6",
   807 => x"50c048f6",
   808 => x"bfcef5c0",
   809 => x"87e1c248",
   810 => x"48c3f0c2",
   811 => x"c27e50c0",
   812 => x"49bff2ef",
   813 => x"bfe2e7c2",
   814 => x"04aa714a",
   815 => x"c287f6fb",
   816 => x"05bfd3f4",
   817 => x"c287c8c0",
   818 => x"02bfeeef",
   819 => x"c287f8c1",
   820 => x"49bfdee7",
   821 => x"7087c9e9",
   822 => x"e2e7c249",
   823 => x"48a6c459",
   824 => x"bfdee7c2",
   825 => x"eeefc278",
   826 => x"d8c002bf",
   827 => x"4966c487",
   828 => x"ffffffcf",
   829 => x"02a999f8",
   830 => x"c087c5c0",
   831 => x"87e1c04c",
   832 => x"dcc04cc1",
   833 => x"4966c487",
   834 => x"99f8ffcf",
   835 => x"c8c002a9",
   836 => x"48a6c887",
   837 => x"c5c078c0",
   838 => x"48a6c887",
   839 => x"66c878c1",
   840 => x"059c744c",
   841 => x"c487e0c0",
   842 => x"89c24966",
   843 => x"bfe6efc2",
   844 => x"f3c2914a",
   845 => x"c24abfff",
   846 => x"7248dae7",
   847 => x"e7c278a1",
   848 => x"78c048e2",
   849 => x"c087def9",
   850 => x"e78ef448",
   851 => x"000087ca",
   852 => x"ffff0000",
   853 => x"0d5effff",
   854 => x"0d670000",
   855 => x"41460000",
   856 => x"20323354",
   857 => x"46002020",
   858 => x"36315441",
   859 => x"00202020",
   860 => x"d8f4c21e",
   861 => x"a8dd48bf",
   862 => x"c087c905",
   863 => x"7087dbfd",
   864 => x"87c84a49",
   865 => x"c348d4ff",
   866 => x"4a6878ff",
   867 => x"4f264872",
   868 => x"d8f4c21e",
   869 => x"a8dd48bf",
   870 => x"c087c605",
   871 => x"d987e7fc",
   872 => x"48d4ff87",
   873 => x"ff78ffc3",
   874 => x"e1c848d0",
   875 => x"48d4ff78",
   876 => x"f4c278d4",
   877 => x"d4ff48d7",
   878 => x"4f2650bf",
   879 => x"48d0ff1e",
   880 => x"2678e0c0",
   881 => x"e7fe1e4f",
   882 => x"99497087",
   883 => x"c087c602",
   884 => x"f105a9fb",
   885 => x"26487187",
   886 => x"5b5e0e4f",
   887 => x"4b710e5c",
   888 => x"cbfe4cc0",
   889 => x"99497087",
   890 => x"87f9c002",
   891 => x"02a9ecc0",
   892 => x"c087f2c0",
   893 => x"c002a9fb",
   894 => x"66cc87eb",
   895 => x"c703acb7",
   896 => x"0266d087",
   897 => x"537187c2",
   898 => x"c2029971",
   899 => x"fd84c187",
   900 => x"497087de",
   901 => x"87cd0299",
   902 => x"02a9ecc0",
   903 => x"fbc087c7",
   904 => x"d5ff05a9",
   905 => x"0266d087",
   906 => x"97c087c3",
   907 => x"a9ecc07b",
   908 => x"7487c405",
   909 => x"7487c54a",
   910 => x"8a0ac04a",
   911 => x"87c24872",
   912 => x"4c264d26",
   913 => x"4f264b26",
   914 => x"87e4fc1e",
   915 => x"f0c04970",
   916 => x"ca04a9b7",
   917 => x"b7f9c087",
   918 => x"87c301a9",
   919 => x"c189f0c0",
   920 => x"04a9b7c1",
   921 => x"dac187ca",
   922 => x"c301a9b7",
   923 => x"89f7c087",
   924 => x"4f264871",
   925 => x"5c5b5e0e",
   926 => x"fc4c710e",
   927 => x"1ec187d2",
   928 => x"741e66d0",
   929 => x"87d1fd49",
   930 => x"4b7086c8",
   931 => x"c087edfc",
   932 => x"c203abb7",
   933 => x"cc8b0b87",
   934 => x"03abb766",
   935 => x"a37487cf",
   936 => x"c083c149",
   937 => x"66cc51e0",
   938 => x"f104abb7",
   939 => x"49a37487",
   940 => x"cdfe51c0",
   941 => x"5b5e0e87",
   942 => x"4a710e5c",
   943 => x"724cd4ff",
   944 => x"87eac049",
   945 => x"029b4b70",
   946 => x"8bc187c2",
   947 => x"c848d0ff",
   948 => x"d5c178c5",
   949 => x"c649737c",
   950 => x"cfe1c231",
   951 => x"484abf97",
   952 => x"7c70b071",
   953 => x"c448d0ff",
   954 => x"fd487378",
   955 => x"5e0e87d4",
   956 => x"0e5d5c5b",
   957 => x"4c7186f4",
   958 => x"c048a6c4",
   959 => x"7ea4c878",
   960 => x"49bf976e",
   961 => x"05a9c1c1",
   962 => x"a4c987dd",
   963 => x"49699749",
   964 => x"05a9d2c1",
   965 => x"a4ca87d1",
   966 => x"49699749",
   967 => x"05a9c3c1",
   968 => x"48df87c5",
   969 => x"f987e1c2",
   970 => x"4bc087e6",
   971 => x"97cdffc0",
   972 => x"a9c049bf",
   973 => x"fa87cf04",
   974 => x"83c187cb",
   975 => x"97cdffc0",
   976 => x"06ab49bf",
   977 => x"ffc087f1",
   978 => x"02bf97cd",
   979 => x"dff887cf",
   980 => x"99497087",
   981 => x"c087c602",
   982 => x"f105a9ec",
   983 => x"f84bc087",
   984 => x"4d7087ce",
   985 => x"cc87c9f8",
   986 => x"c3f858a6",
   987 => x"c14a7087",
   988 => x"bf976e83",
   989 => x"c702ad49",
   990 => x"adffc087",
   991 => x"87eac005",
   992 => x"9749a4c9",
   993 => x"66c84969",
   994 => x"87c702a9",
   995 => x"a8ffc048",
   996 => x"ca87d705",
   997 => x"699749a4",
   998 => x"c602aa49",
   999 => x"aaffc087",
  1000 => x"c487c705",
  1001 => x"78c148a6",
  1002 => x"ecc087d3",
  1003 => x"87c602ad",
  1004 => x"05adfbc0",
  1005 => x"4bc087c7",
  1006 => x"c148a6c4",
  1007 => x"0266c478",
  1008 => x"f787dcfe",
  1009 => x"487387f6",
  1010 => x"f3f98ef4",
  1011 => x"5e0e0087",
  1012 => x"0e5d5c5b",
  1013 => x"c04b711e",
  1014 => x"04ab4d4c",
  1015 => x"c087e8c0",
  1016 => x"751eeefb",
  1017 => x"87c4029d",
  1018 => x"87c24ac0",
  1019 => x"49724ac1",
  1020 => x"c487c3ee",
  1021 => x"c17e7086",
  1022 => x"c2056e84",
  1023 => x"c14c7387",
  1024 => x"06ac7385",
  1025 => x"6e87d8ff",
  1026 => x"4d262648",
  1027 => x"4b264c26",
  1028 => x"5e0e4f26",
  1029 => x"0e5d5c5b",
  1030 => x"494c711e",
  1031 => x"f4c291de",
  1032 => x"85714df1",
  1033 => x"c1026d97",
  1034 => x"f4c287dd",
  1035 => x"744abfdc",
  1036 => x"fe497282",
  1037 => x"7e7087d8",
  1038 => x"f3c0026e",
  1039 => x"e4f4c287",
  1040 => x"cb4a6e4b",
  1041 => x"dfc1ff49",
  1042 => x"cb4b7487",
  1043 => x"d8e2c193",
  1044 => x"c183c483",
  1045 => x"747bcbc2",
  1046 => x"c8cbc149",
  1047 => x"c27b7587",
  1048 => x"bf97f0f4",
  1049 => x"f4c21e49",
  1050 => x"dfc149e4",
  1051 => x"86c487d2",
  1052 => x"cac14974",
  1053 => x"49c087ef",
  1054 => x"87ceccc1",
  1055 => x"48d8f4c2",
  1056 => x"49c178c0",
  1057 => x"2687c3dd",
  1058 => x"4c87fffd",
  1059 => x"6964616f",
  1060 => x"2e2e676e",
  1061 => x"5e0e002e",
  1062 => x"710e5c5b",
  1063 => x"f4c24a4b",
  1064 => x"7282bfdc",
  1065 => x"87e6fc49",
  1066 => x"029c4c70",
  1067 => x"ea4987c4",
  1068 => x"f4c287cc",
  1069 => x"78c048dc",
  1070 => x"cddc49c1",
  1071 => x"87ccfd87",
  1072 => x"5c5b5e0e",
  1073 => x"86f40e5d",
  1074 => x"4de6e7c2",
  1075 => x"a6c44cc0",
  1076 => x"c278c048",
  1077 => x"49bfdcf4",
  1078 => x"c106a9c0",
  1079 => x"e7c287c1",
  1080 => x"029848e6",
  1081 => x"c087f8c0",
  1082 => x"c81eeefb",
  1083 => x"87c70266",
  1084 => x"c048a6c4",
  1085 => x"c487c578",
  1086 => x"78c148a6",
  1087 => x"e94966c4",
  1088 => x"86c487f4",
  1089 => x"84c14d70",
  1090 => x"c14866c4",
  1091 => x"58a6c880",
  1092 => x"bfdcf4c2",
  1093 => x"c603ac49",
  1094 => x"059d7587",
  1095 => x"c087c8ff",
  1096 => x"029d754c",
  1097 => x"c087e0c3",
  1098 => x"c81eeefb",
  1099 => x"87c70266",
  1100 => x"c048a6cc",
  1101 => x"cc87c578",
  1102 => x"78c148a6",
  1103 => x"e84966cc",
  1104 => x"86c487f4",
  1105 => x"026e7e70",
  1106 => x"6e87e9c2",
  1107 => x"9781cb49",
  1108 => x"99d04969",
  1109 => x"87d6c102",
  1110 => x"4ad6c2c1",
  1111 => x"91cb4974",
  1112 => x"81d8e2c1",
  1113 => x"81c87972",
  1114 => x"7451ffc3",
  1115 => x"c291de49",
  1116 => x"714df1f4",
  1117 => x"97c1c285",
  1118 => x"49a5c17d",
  1119 => x"c251e0c0",
  1120 => x"bf97f6ef",
  1121 => x"c187d202",
  1122 => x"4ba5c284",
  1123 => x"4af6efc2",
  1124 => x"fcfe49db",
  1125 => x"dbc187d2",
  1126 => x"49a5cd87",
  1127 => x"84c151c0",
  1128 => x"6e4ba5c2",
  1129 => x"fe49cb4a",
  1130 => x"c187fdfb",
  1131 => x"c0c187c6",
  1132 => x"49744ad2",
  1133 => x"e2c191cb",
  1134 => x"797281d8",
  1135 => x"97f6efc2",
  1136 => x"87d802bf",
  1137 => x"91de4974",
  1138 => x"f4c284c1",
  1139 => x"83714bf1",
  1140 => x"4af6efc2",
  1141 => x"fbfe49dd",
  1142 => x"87d887ce",
  1143 => x"93de4b74",
  1144 => x"83f1f4c2",
  1145 => x"c049a3cb",
  1146 => x"7384c151",
  1147 => x"49cb4a6e",
  1148 => x"87f4fafe",
  1149 => x"c14866c4",
  1150 => x"58a6c880",
  1151 => x"c003acc7",
  1152 => x"056e87c5",
  1153 => x"7487e0fc",
  1154 => x"f78ef448",
  1155 => x"731e87fc",
  1156 => x"494b711e",
  1157 => x"e2c191cb",
  1158 => x"a1c881d8",
  1159 => x"cfe1c24a",
  1160 => x"c9501248",
  1161 => x"ffc04aa1",
  1162 => x"501248cd",
  1163 => x"f4c281ca",
  1164 => x"501148f0",
  1165 => x"97f0f4c2",
  1166 => x"c01e49bf",
  1167 => x"ffd7c149",
  1168 => x"d8f4c287",
  1169 => x"c178de48",
  1170 => x"87fed549",
  1171 => x"87fef626",
  1172 => x"494a711e",
  1173 => x"e2c191cb",
  1174 => x"81c881d8",
  1175 => x"f4c24811",
  1176 => x"f4c258dc",
  1177 => x"78c048dc",
  1178 => x"ddd549c1",
  1179 => x"1e4f2687",
  1180 => x"c4c149c0",
  1181 => x"4f2687d4",
  1182 => x"0299711e",
  1183 => x"e3c187d2",
  1184 => x"50c048ed",
  1185 => x"c9c180f7",
  1186 => x"e2c140d0",
  1187 => x"87ce78d1",
  1188 => x"48e9e3c1",
  1189 => x"78cae2c1",
  1190 => x"c9c180fc",
  1191 => x"4f2678ef",
  1192 => x"5c5b5e0e",
  1193 => x"4a4c710e",
  1194 => x"e2c192cb",
  1195 => x"a2c882d8",
  1196 => x"4ba2c949",
  1197 => x"1e4b6b97",
  1198 => x"1e496997",
  1199 => x"491282ca",
  1200 => x"87f5e4c0",
  1201 => x"c1d449c0",
  1202 => x"c1497487",
  1203 => x"f887d6c1",
  1204 => x"87f8f48e",
  1205 => x"711e731e",
  1206 => x"c3ff494b",
  1207 => x"fe497387",
  1208 => x"e9f487fe",
  1209 => x"1e731e87",
  1210 => x"a3c64b71",
  1211 => x"87db024a",
  1212 => x"d6028ac1",
  1213 => x"c1028a87",
  1214 => x"028a87da",
  1215 => x"8a87fcc0",
  1216 => x"87e1c002",
  1217 => x"87cb028a",
  1218 => x"c787dbc1",
  1219 => x"87c0fd49",
  1220 => x"c287dec1",
  1221 => x"02bfdcf4",
  1222 => x"4887cbc1",
  1223 => x"f4c288c1",
  1224 => x"c1c158e0",
  1225 => x"e0f4c287",
  1226 => x"f9c002bf",
  1227 => x"dcf4c287",
  1228 => x"80c148bf",
  1229 => x"58e0f4c2",
  1230 => x"c287ebc0",
  1231 => x"49bfdcf4",
  1232 => x"f4c289c6",
  1233 => x"b7c059e0",
  1234 => x"87da03a9",
  1235 => x"48dcf4c2",
  1236 => x"87d278c0",
  1237 => x"bfe0f4c2",
  1238 => x"c287cb02",
  1239 => x"48bfdcf4",
  1240 => x"f4c280c6",
  1241 => x"49c058e0",
  1242 => x"7387dfd1",
  1243 => x"f4fec049",
  1244 => x"87daf287",
  1245 => x"711e731e",
  1246 => x"d8f4c24b",
  1247 => x"c078dd48",
  1248 => x"87c6d149",
  1249 => x"fec04973",
  1250 => x"c1f287db",
  1251 => x"5b5e0e87",
  1252 => x"4c710e5c",
  1253 => x"741e66cc",
  1254 => x"c193cb4b",
  1255 => x"c483d8e2",
  1256 => x"496a4aa3",
  1257 => x"87d0f4fe",
  1258 => x"7bcec8c1",
  1259 => x"d449a3c8",
  1260 => x"a3c95166",
  1261 => x"5166d849",
  1262 => x"dc49a3ca",
  1263 => x"f1265166",
  1264 => x"5e0e87ca",
  1265 => x"0e5d5c5b",
  1266 => x"dc86ccff",
  1267 => x"a6c859a6",
  1268 => x"c478c048",
  1269 => x"66c8c180",
  1270 => x"c180c478",
  1271 => x"c180c478",
  1272 => x"e0f4c278",
  1273 => x"c278c148",
  1274 => x"48bfd8f4",
  1275 => x"cb05a8de",
  1276 => x"87ccf387",
  1277 => x"a6cc4970",
  1278 => x"87cace59",
  1279 => x"e787d1e6",
  1280 => x"ebe587c3",
  1281 => x"c04c7087",
  1282 => x"c102acfb",
  1283 => x"66d887d8",
  1284 => x"87cac105",
  1285 => x"c11e1ec0",
  1286 => x"fbe3c11e",
  1287 => x"fd49c01e",
  1288 => x"86d087eb",
  1289 => x"02acfbc0",
  1290 => x"c4c187d9",
  1291 => x"82c44a66",
  1292 => x"81c7496a",
  1293 => x"1ec15174",
  1294 => x"496a1ed8",
  1295 => x"d8e681c8",
  1296 => x"c186c887",
  1297 => x"c04866c8",
  1298 => x"87c701a8",
  1299 => x"c148a6c8",
  1300 => x"c187ce78",
  1301 => x"c14866c8",
  1302 => x"58a6d088",
  1303 => x"e4e587c3",
  1304 => x"48a6d087",
  1305 => x"9c7478c2",
  1306 => x"87d6cc02",
  1307 => x"c14866c8",
  1308 => x"03a866cc",
  1309 => x"c487cbcc",
  1310 => x"78c048a6",
  1311 => x"78c080d8",
  1312 => x"7087ede3",
  1313 => x"4866d84c",
  1314 => x"c605a8dd",
  1315 => x"48a6dc87",
  1316 => x"c17866d8",
  1317 => x"c005acd0",
  1318 => x"d3e387e8",
  1319 => x"87d0e387",
  1320 => x"ecc04c70",
  1321 => x"87c505ac",
  1322 => x"7087dae4",
  1323 => x"acd0c14c",
  1324 => x"d487c805",
  1325 => x"80c14866",
  1326 => x"c158a6d8",
  1327 => x"ff02acd0",
  1328 => x"e0c087d8",
  1329 => x"66d848a6",
  1330 => x"4866dc78",
  1331 => x"a866e0c0",
  1332 => x"87c0ca05",
  1333 => x"48a6e4c0",
  1334 => x"80c478c0",
  1335 => x"4d7478c0",
  1336 => x"028dfbc0",
  1337 => x"c987c6c9",
  1338 => x"87db028d",
  1339 => x"c1028dc2",
  1340 => x"8dc987f4",
  1341 => x"87cbc402",
  1342 => x"c1028dc4",
  1343 => x"8dc187c1",
  1344 => x"87ffc302",
  1345 => x"c887e0c8",
  1346 => x"91cb4966",
  1347 => x"8166c4c1",
  1348 => x"6a4aa1c4",
  1349 => x"c11e717e",
  1350 => x"c448fdde",
  1351 => x"a1cc4966",
  1352 => x"7141204a",
  1353 => x"f8ff05aa",
  1354 => x"26511087",
  1355 => x"f4cdc149",
  1356 => x"87d1e279",
  1357 => x"e8c04c70",
  1358 => x"78c148a6",
  1359 => x"c487eec7",
  1360 => x"f0c048a6",
  1361 => x"87e8e078",
  1362 => x"ecc04c70",
  1363 => x"c3c002ac",
  1364 => x"5ca6c887",
  1365 => x"02acecc0",
  1366 => x"d3e087cc",
  1367 => x"c04c7087",
  1368 => x"ff05acec",
  1369 => x"ecc087f4",
  1370 => x"c3c002ac",
  1371 => x"87c0e087",
  1372 => x"d81e66c4",
  1373 => x"d81e4966",
  1374 => x"c11e4966",
  1375 => x"d81efbe3",
  1376 => x"c8f84966",
  1377 => x"ca1ec087",
  1378 => x"66e0c01e",
  1379 => x"c191cb49",
  1380 => x"d88166dc",
  1381 => x"a1c448a6",
  1382 => x"bf66d878",
  1383 => x"87f9e049",
  1384 => x"b7c086d8",
  1385 => x"cac106a8",
  1386 => x"de1ec187",
  1387 => x"bf66c81e",
  1388 => x"87e5e049",
  1389 => x"497086c8",
  1390 => x"8808c048",
  1391 => x"58a6ecc0",
  1392 => x"06a8b7c0",
  1393 => x"c087ecc0",
  1394 => x"dd4866e8",
  1395 => x"c003a8b7",
  1396 => x"bf6e87e1",
  1397 => x"66e8c049",
  1398 => x"51e0c081",
  1399 => x"4966e8c0",
  1400 => x"bf6e81c1",
  1401 => x"51c1c281",
  1402 => x"4966e8c0",
  1403 => x"bf6e81c2",
  1404 => x"d051c081",
  1405 => x"80c14866",
  1406 => x"4858a6d4",
  1407 => x"78c180d8",
  1408 => x"e187eac4",
  1409 => x"ecc087c2",
  1410 => x"fbe058a6",
  1411 => x"a6f0c087",
  1412 => x"a8ecc058",
  1413 => x"87c9c005",
  1414 => x"e8c048a6",
  1415 => x"c4c07866",
  1416 => x"cbddff87",
  1417 => x"4966c887",
  1418 => x"c4c191cb",
  1419 => x"80714866",
  1420 => x"c458a6c8",
  1421 => x"82c84a66",
  1422 => x"ca4966c4",
  1423 => x"66e8c081",
  1424 => x"66ecc051",
  1425 => x"c081c149",
  1426 => x"c18966e8",
  1427 => x"70307148",
  1428 => x"7189c149",
  1429 => x"f8c27a97",
  1430 => x"c049bfcd",
  1431 => x"972966e8",
  1432 => x"71484a6a",
  1433 => x"a6f4c098",
  1434 => x"4966c458",
  1435 => x"7e6981c4",
  1436 => x"4866e0c0",
  1437 => x"02a866dc",
  1438 => x"dc87c8c0",
  1439 => x"78c048a6",
  1440 => x"dc87c5c0",
  1441 => x"78c148a6",
  1442 => x"c01e66dc",
  1443 => x"66c81ee0",
  1444 => x"c4ddff49",
  1445 => x"7086c887",
  1446 => x"acb7c04c",
  1447 => x"87d6c106",
  1448 => x"8074486e",
  1449 => x"e0c07e70",
  1450 => x"6e897449",
  1451 => x"fadec14b",
  1452 => x"e7fe714a",
  1453 => x"486e87f2",
  1454 => x"7e7080c2",
  1455 => x"4866e4c0",
  1456 => x"e8c080c1",
  1457 => x"f0c058a6",
  1458 => x"81c14966",
  1459 => x"c002a970",
  1460 => x"4dc087c5",
  1461 => x"c187c2c0",
  1462 => x"c21e754d",
  1463 => x"e0c049a4",
  1464 => x"70887148",
  1465 => x"66c81e49",
  1466 => x"ecdbff49",
  1467 => x"c086c887",
  1468 => x"ff01a8b7",
  1469 => x"e4c087c6",
  1470 => x"d3c00266",
  1471 => x"4966c487",
  1472 => x"e4c081c9",
  1473 => x"66c45166",
  1474 => x"e0cac148",
  1475 => x"87cec078",
  1476 => x"c94966c4",
  1477 => x"c451c281",
  1478 => x"cbc14866",
  1479 => x"e8c078d4",
  1480 => x"78c148a6",
  1481 => x"ff87c6c0",
  1482 => x"7087dada",
  1483 => x"66e8c04c",
  1484 => x"87f5c002",
  1485 => x"cc4866c8",
  1486 => x"c004a866",
  1487 => x"66c887cb",
  1488 => x"cc80c148",
  1489 => x"e0c058a6",
  1490 => x"4866cc87",
  1491 => x"a6d088c1",
  1492 => x"87d5c058",
  1493 => x"05acc6c1",
  1494 => x"d087c8c0",
  1495 => x"80c14866",
  1496 => x"ff58a6d4",
  1497 => x"7087ded9",
  1498 => x"4866d44c",
  1499 => x"a6d880c1",
  1500 => x"029c7458",
  1501 => x"c887cbc0",
  1502 => x"ccc14866",
  1503 => x"f304a866",
  1504 => x"d8ff87f5",
  1505 => x"66c887f6",
  1506 => x"03a8c748",
  1507 => x"c287e5c0",
  1508 => x"c048e0f4",
  1509 => x"4966c878",
  1510 => x"c4c191cb",
  1511 => x"a1c48166",
  1512 => x"c04a6a4a",
  1513 => x"66c87952",
  1514 => x"cc80c148",
  1515 => x"a8c758a6",
  1516 => x"87dbff04",
  1517 => x"e18eccff",
  1518 => x"203a87d0",
  1519 => x"50494400",
  1520 => x"69775320",
  1521 => x"65686374",
  1522 => x"731e0073",
  1523 => x"9b4b711e",
  1524 => x"c287c602",
  1525 => x"c048dcf4",
  1526 => x"c21ec778",
  1527 => x"49bfdcf4",
  1528 => x"d8e2c11e",
  1529 => x"d8f4c21e",
  1530 => x"d5ef49bf",
  1531 => x"c286cc87",
  1532 => x"49bfd8f4",
  1533 => x"7387c1ea",
  1534 => x"87c8029b",
  1535 => x"49d8e2c1",
  1536 => x"87f3edc0",
  1537 => x"1e87c7e0",
  1538 => x"c187cfc7",
  1539 => x"87fafe49",
  1540 => x"87efeafe",
  1541 => x"cd029870",
  1542 => x"c8f2fe87",
  1543 => x"02987087",
  1544 => x"4ac187c4",
  1545 => x"4ac087c2",
  1546 => x"ce059a72",
  1547 => x"c11ec087",
  1548 => x"c049dce1",
  1549 => x"c487def9",
  1550 => x"c187fe86",
  1551 => x"c087fac0",
  1552 => x"e7e1c11e",
  1553 => x"ccf9c049",
  1554 => x"c11ec087",
  1555 => x"7087c0c3",
  1556 => x"c0f9c049",
  1557 => x"87c1c387",
  1558 => x"4f268ef8",
  1559 => x"66204453",
  1560 => x"656c6961",
  1561 => x"42002e64",
  1562 => x"69746f6f",
  1563 => x"2e2e676e",
  1564 => x"c21e002e",
  1565 => x"c048dcf4",
  1566 => x"d8f4c278",
  1567 => x"fe78c048",
  1568 => x"c4c187c5",
  1569 => x"48c087e6",
  1570 => x"20804f26",
  1571 => x"74697845",
  1572 => x"42208000",
  1573 => x"006b6361",
  1574 => x"00001250",
  1575 => x"00002d31",
  1576 => x"50000000",
  1577 => x"4f000012",
  1578 => x"0000002d",
  1579 => x"12500000",
  1580 => x"2d6d0000",
  1581 => x"00000000",
  1582 => x"00125000",
  1583 => x"002d8b00",
  1584 => x"00000000",
  1585 => x"00001250",
  1586 => x"00002da9",
  1587 => x"50000000",
  1588 => x"c7000012",
  1589 => x"0000002d",
  1590 => x"12500000",
  1591 => x"2de50000",
  1592 => x"00000000",
  1593 => x"00125000",
  1594 => x"00000000",
  1595 => x"00000000",
  1596 => x"000012e5",
  1597 => x"00000000",
  1598 => x"4c000000",
  1599 => x"2064616f",
  1600 => x"1e002e2a",
  1601 => x"c048f0fe",
  1602 => x"7909cd78",
  1603 => x"1e4f2609",
  1604 => x"bff0fe1e",
  1605 => x"2626487e",
  1606 => x"f0fe1e4f",
  1607 => x"2678c148",
  1608 => x"f0fe1e4f",
  1609 => x"2678c048",
  1610 => x"4a711e4f",
  1611 => x"265252c0",
  1612 => x"5b5e0e4f",
  1613 => x"f40e5d5c",
  1614 => x"974d7186",
  1615 => x"a5c17e6d",
  1616 => x"486c974c",
  1617 => x"6e58a6c8",
  1618 => x"a866c448",
  1619 => x"ff87c505",
  1620 => x"87e6c048",
  1621 => x"c287caff",
  1622 => x"6c9749a5",
  1623 => x"4ba3714b",
  1624 => x"974b6b97",
  1625 => x"486e7e6c",
  1626 => x"a6c880c1",
  1627 => x"cc98c758",
  1628 => x"977058a6",
  1629 => x"87e1fe7c",
  1630 => x"8ef44873",
  1631 => x"4c264d26",
  1632 => x"4f264b26",
  1633 => x"5c5b5e0e",
  1634 => x"7186f40e",
  1635 => x"4a66d84c",
  1636 => x"c29affc3",
  1637 => x"6c974ba4",
  1638 => x"49a17349",
  1639 => x"6c975172",
  1640 => x"c1486e7e",
  1641 => x"58a6c880",
  1642 => x"a6cc98c7",
  1643 => x"f4547058",
  1644 => x"87caff8e",
  1645 => x"e8fd1e1e",
  1646 => x"4abfe087",
  1647 => x"c0e0c049",
  1648 => x"87cb0299",
  1649 => x"f8c21e72",
  1650 => x"f7fe49c3",
  1651 => x"fc86c487",
  1652 => x"7e7087fd",
  1653 => x"2687c2fd",
  1654 => x"c21e4f26",
  1655 => x"fd49c3f8",
  1656 => x"e6c187c7",
  1657 => x"dafc49f4",
  1658 => x"87c8c487",
  1659 => x"ff1e4f26",
  1660 => x"e1c848d0",
  1661 => x"48d4ff78",
  1662 => x"66c478c5",
  1663 => x"c387c302",
  1664 => x"66c878e0",
  1665 => x"ff87c602",
  1666 => x"f0c348d4",
  1667 => x"48d4ff78",
  1668 => x"d0ff7871",
  1669 => x"78e1c848",
  1670 => x"2678e0c0",
  1671 => x"5b5e0e4f",
  1672 => x"4c710e5c",
  1673 => x"49c3f8c2",
  1674 => x"7087c6fc",
  1675 => x"aab7c04a",
  1676 => x"87e3c204",
  1677 => x"05aae0c3",
  1678 => x"ebc187c9",
  1679 => x"78c148e7",
  1680 => x"c387d4c2",
  1681 => x"c905aaf0",
  1682 => x"e3ebc187",
  1683 => x"c178c148",
  1684 => x"ebc187f5",
  1685 => x"c702bfe7",
  1686 => x"c24b7287",
  1687 => x"87c2b3c0",
  1688 => x"9c744b72",
  1689 => x"c187d105",
  1690 => x"1ebfe3eb",
  1691 => x"bfe7ebc1",
  1692 => x"fd49721e",
  1693 => x"86c887f8",
  1694 => x"bfe3ebc1",
  1695 => x"87e0c002",
  1696 => x"b7c44973",
  1697 => x"edc19129",
  1698 => x"4a7381c3",
  1699 => x"92c29acf",
  1700 => x"307248c1",
  1701 => x"baff4a70",
  1702 => x"98694872",
  1703 => x"87db7970",
  1704 => x"b7c44973",
  1705 => x"edc19129",
  1706 => x"4a7381c3",
  1707 => x"92c29acf",
  1708 => x"307248c3",
  1709 => x"69484a70",
  1710 => x"c17970b0",
  1711 => x"c048e7eb",
  1712 => x"e3ebc178",
  1713 => x"c278c048",
  1714 => x"f949c3f8",
  1715 => x"4a7087e3",
  1716 => x"03aab7c0",
  1717 => x"c087ddfd",
  1718 => x"2687c248",
  1719 => x"264c264d",
  1720 => x"004f264b",
  1721 => x"00000000",
  1722 => x"1e000000",
  1723 => x"fc494a71",
  1724 => x"4f2687eb",
  1725 => x"724ac01e",
  1726 => x"c191c449",
  1727 => x"c081c3ed",
  1728 => x"d082c179",
  1729 => x"ee04aab7",
  1730 => x"0e4f2687",
  1731 => x"5d5c5b5e",
  1732 => x"f84d710e",
  1733 => x"4a7587cb",
  1734 => x"922ab7c4",
  1735 => x"82c3edc1",
  1736 => x"9ccf4c75",
  1737 => x"496a94c2",
  1738 => x"c32b744b",
  1739 => x"7448c29b",
  1740 => x"ff4c7030",
  1741 => x"714874bc",
  1742 => x"f77a7098",
  1743 => x"487387db",
  1744 => x"0087d8fe",
  1745 => x"00000000",
  1746 => x"00000000",
  1747 => x"00000000",
  1748 => x"00000000",
  1749 => x"00000000",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"00000000",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"1e000000",
  1761 => x"c848d0ff",
  1762 => x"487178e1",
  1763 => x"7808d4ff",
  1764 => x"ff4866c4",
  1765 => x"267808d4",
  1766 => x"4a711e4f",
  1767 => x"1e4966c4",
  1768 => x"deff4972",
  1769 => x"48d0ff87",
  1770 => x"2678e0c0",
  1771 => x"731e4f26",
  1772 => x"c84b711e",
  1773 => x"731e4966",
  1774 => x"a2e0c14a",
  1775 => x"87d9ff49",
  1776 => x"2687c426",
  1777 => x"264c264d",
  1778 => x"1e4f264b",
  1779 => x"c34ad4ff",
  1780 => x"d0ff7aff",
  1781 => x"78e1c848",
  1782 => x"f8c27ade",
  1783 => x"497abfcd",
  1784 => x"7028c848",
  1785 => x"d048717a",
  1786 => x"717a7028",
  1787 => x"7028d848",
  1788 => x"48d0ff7a",
  1789 => x"2678e0c0",
  1790 => x"5b5e0e4f",
  1791 => x"710e5d5c",
  1792 => x"cdf8c24c",
  1793 => x"744b4dbf",
  1794 => x"9b66d02b",
  1795 => x"66d483c1",
  1796 => x"87c204ab",
  1797 => x"4a744bc0",
  1798 => x"724966d0",
  1799 => x"75b9ff31",
  1800 => x"72487399",
  1801 => x"484a7030",
  1802 => x"f8c2b071",
  1803 => x"dafe58d1",
  1804 => x"264d2687",
  1805 => x"264b264c",
  1806 => x"5b5e0e4f",
  1807 => x"1e0e5d5c",
  1808 => x"f8c24c71",
  1809 => x"4ac04bd1",
  1810 => x"fe49f4c0",
  1811 => x"7487f6d1",
  1812 => x"d1f8c21e",
  1813 => x"d8eefe49",
  1814 => x"7086c487",
  1815 => x"eac00298",
  1816 => x"a61ec487",
  1817 => x"f8c21e4d",
  1818 => x"f4fe49d1",
  1819 => x"86c887c6",
  1820 => x"d6029870",
  1821 => x"c14a7587",
  1822 => x"c449c1f3",
  1823 => x"e9cffe4b",
  1824 => x"02987087",
  1825 => x"48c087ca",
  1826 => x"c087edc0",
  1827 => x"87e8c048",
  1828 => x"c187f3c0",
  1829 => x"987087c4",
  1830 => x"c087c802",
  1831 => x"987087fc",
  1832 => x"c287f805",
  1833 => x"02bff1f8",
  1834 => x"f8c287cc",
  1835 => x"f8c248cd",
  1836 => x"fc78bff1",
  1837 => x"48c187d5",
  1838 => x"264d2626",
  1839 => x"264b264c",
  1840 => x"52415b4f",
  1841 => x"c01e0043",
  1842 => x"d1f8c21e",
  1843 => x"fcf0fe49",
  1844 => x"e9f8c287",
  1845 => x"2678c048",
  1846 => x"5e0e4f26",
  1847 => x"0e5d5c5b",
  1848 => x"a6c486f4",
  1849 => x"c278c048",
  1850 => x"48bfe9f8",
  1851 => x"03a8b7c3",
  1852 => x"f8c287d1",
  1853 => x"c148bfe9",
  1854 => x"edf8c280",
  1855 => x"48fbc058",
  1856 => x"c287e2c6",
  1857 => x"fe49d1f8",
  1858 => x"7087fdf5",
  1859 => x"e9f8c24c",
  1860 => x"8ac34abf",
  1861 => x"c187d802",
  1862 => x"cbc5028a",
  1863 => x"c2028a87",
  1864 => x"028a87f6",
  1865 => x"8a87cdc1",
  1866 => x"87e2c302",
  1867 => x"c087e1c5",
  1868 => x"c44a754d",
  1869 => x"c3fbc192",
  1870 => x"e5f8c282",
  1871 => x"70807548",
  1872 => x"bf976e7e",
  1873 => x"6e4b494b",
  1874 => x"50a3c148",
  1875 => x"4811816a",
  1876 => x"7058a6cc",
  1877 => x"87c402ac",
  1878 => x"50c0486e",
  1879 => x"c70566c8",
  1880 => x"e9f8c287",
  1881 => x"78a5c448",
  1882 => x"b7c485c1",
  1883 => x"c0ff04ad",
  1884 => x"87dcc487",
  1885 => x"bff5f8c2",
  1886 => x"a8b7c848",
  1887 => x"ca87d101",
  1888 => x"87cc02ac",
  1889 => x"c702accd",
  1890 => x"acb7c087",
  1891 => x"87f3c003",
  1892 => x"bff5f8c2",
  1893 => x"abb7c84b",
  1894 => x"c287d203",
  1895 => x"7349f9f8",
  1896 => x"51e0c081",
  1897 => x"b7c883c1",
  1898 => x"eeff04ab",
  1899 => x"c1f9c287",
  1900 => x"50d2c148",
  1901 => x"c150cfc1",
  1902 => x"50c050cd",
  1903 => x"78c380e4",
  1904 => x"c287cdc3",
  1905 => x"49bff5f8",
  1906 => x"c280c148",
  1907 => x"4858f9f8",
  1908 => x"7481a0c4",
  1909 => x"87f8c251",
  1910 => x"acb7f0c0",
  1911 => x"c087da04",
  1912 => x"01acb7f9",
  1913 => x"f8c287d3",
  1914 => x"ca49bfed",
  1915 => x"c04a7491",
  1916 => x"f8c28af0",
  1917 => x"a17248ed",
  1918 => x"02acca78",
  1919 => x"cd87c6c0",
  1920 => x"cbc205ac",
  1921 => x"e9f8c287",
  1922 => x"c278c348",
  1923 => x"f0c087c2",
  1924 => x"db04acb7",
  1925 => x"b7f9c087",
  1926 => x"d3c001ac",
  1927 => x"f1f8c287",
  1928 => x"91d049bf",
  1929 => x"f0c04a74",
  1930 => x"f1f8c28a",
  1931 => x"78a17248",
  1932 => x"acb7c1c1",
  1933 => x"87dbc004",
  1934 => x"acb7c6c1",
  1935 => x"87d3c001",
  1936 => x"bff1f8c2",
  1937 => x"7491d049",
  1938 => x"8af7c04a",
  1939 => x"48f1f8c2",
  1940 => x"ca78a172",
  1941 => x"c6c002ac",
  1942 => x"05accd87",
  1943 => x"c287f1c0",
  1944 => x"c348e9f8",
  1945 => x"87e8c078",
  1946 => x"05ace2c0",
  1947 => x"c487c9c0",
  1948 => x"fbc048a6",
  1949 => x"87d8c078",
  1950 => x"c002acca",
  1951 => x"accd87c6",
  1952 => x"87c9c005",
  1953 => x"48e9f8c2",
  1954 => x"c3c078c3",
  1955 => x"5ca6c887",
  1956 => x"03acb7c0",
  1957 => x"4887c4c0",
  1958 => x"c487cac0",
  1959 => x"c6f90266",
  1960 => x"ffc34887",
  1961 => x"f88ef499",
  1962 => x"4f4387cf",
  1963 => x"003d464e",
  1964 => x"00444f4d",
  1965 => x"454d414e",
  1966 => x"46454400",
  1967 => x"544c5541",
  1968 => x"aa00303d",
  1969 => x"b000001e",
  1970 => x"b400001e",
  1971 => x"b900001e",
  1972 => x"1e00001e",
  1973 => x"c848d0ff",
  1974 => x"487178c9",
  1975 => x"7808d4ff",
  1976 => x"711e4f26",
  1977 => x"87eb494a",
  1978 => x"c848d0ff",
  1979 => x"1e4f2678",
  1980 => x"4b711e73",
  1981 => x"bfd1f9c2",
  1982 => x"c287c302",
  1983 => x"d0ff87eb",
  1984 => x"78c9c848",
  1985 => x"e0c04973",
  1986 => x"48d4ffb1",
  1987 => x"f9c27871",
  1988 => x"78c048c5",
  1989 => x"c50266c8",
  1990 => x"49ffc387",
  1991 => x"49c087c2",
  1992 => x"59cdf9c2",
  1993 => x"c60266cc",
  1994 => x"d5d5c587",
  1995 => x"cf87c44a",
  1996 => x"c24affff",
  1997 => x"c25ad1f9",
  1998 => x"c148d1f9",
  1999 => x"2687c478",
  2000 => x"264c264d",
  2001 => x"0e4f264b",
  2002 => x"5d5c5b5e",
  2003 => x"c24a710e",
  2004 => x"4cbfcdf9",
  2005 => x"cb029a72",
  2006 => x"91c84987",
  2007 => x"4be5fbc1",
  2008 => x"87c48371",
  2009 => x"4be5ffc1",
  2010 => x"49134dc0",
  2011 => x"f9c29974",
  2012 => x"ffb9bfc9",
  2013 => x"787148d4",
  2014 => x"852cb7c1",
  2015 => x"04adb7c8",
  2016 => x"f9c287e8",
  2017 => x"c848bfc5",
  2018 => x"c9f9c280",
  2019 => x"87effe58",
  2020 => x"711e731e",
  2021 => x"9a4a134b",
  2022 => x"7287cb02",
  2023 => x"87e7fe49",
  2024 => x"059a4a13",
  2025 => x"dafe87f5",
  2026 => x"f9c21e87",
  2027 => x"c249bfc5",
  2028 => x"c148c5f9",
  2029 => x"c0c478a1",
  2030 => x"db03a9b7",
  2031 => x"48d4ff87",
  2032 => x"bfc9f9c2",
  2033 => x"c5f9c278",
  2034 => x"f9c249bf",
  2035 => x"a1c148c5",
  2036 => x"b7c0c478",
  2037 => x"87e504a9",
  2038 => x"c848d0ff",
  2039 => x"d1f9c278",
  2040 => x"2678c048",
  2041 => x"0000004f",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00005f5f",
  2045 => x"03030000",
  2046 => x"00030300",
  2047 => x"7f7f1400",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
