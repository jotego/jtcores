library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"147f7f14",
     1 => x"2e240000",
     2 => x"123a6b6b",
     3 => x"366a4c00",
     4 => x"32566c18",
     5 => x"4f7e3000",
     6 => x"683a7759",
     7 => x"04000040",
     8 => x"00000307",
     9 => x"1c000000",
    10 => x"0041633e",
    11 => x"41000000",
    12 => x"001c3e63",
    13 => x"3e2a0800",
    14 => x"2a3e1c1c",
    15 => x"08080008",
    16 => x"08083e3e",
    17 => x"80000000",
    18 => x"000060e0",
    19 => x"08080000",
    20 => x"08080808",
    21 => x"00000000",
    22 => x"00006060",
    23 => x"30604000",
    24 => x"03060c18",
    25 => x"7f3e0001",
    26 => x"3e7f4d59",
    27 => x"06040000",
    28 => x"00007f7f",
    29 => x"63420000",
    30 => x"464f5971",
    31 => x"63220000",
    32 => x"367f4949",
    33 => x"161c1800",
    34 => x"107f7f13",
    35 => x"67270000",
    36 => x"397d4545",
    37 => x"7e3c0000",
    38 => x"3079494b",
    39 => x"01010000",
    40 => x"070f7971",
    41 => x"7f360000",
    42 => x"367f4949",
    43 => x"4f060000",
    44 => x"1e3f6949",
    45 => x"00000000",
    46 => x"00006666",
    47 => x"80000000",
    48 => x"000066e6",
    49 => x"08080000",
    50 => x"22221414",
    51 => x"14140000",
    52 => x"14141414",
    53 => x"22220000",
    54 => x"08081414",
    55 => x"03020000",
    56 => x"060f5951",
    57 => x"417f3e00",
    58 => x"1e1f555d",
    59 => x"7f7e0000",
    60 => x"7e7f0909",
    61 => x"7f7f0000",
    62 => x"367f4949",
    63 => x"3e1c0000",
    64 => x"41414163",
    65 => x"7f7f0000",
    66 => x"1c3e6341",
    67 => x"7f7f0000",
    68 => x"41414949",
    69 => x"7f7f0000",
    70 => x"01010909",
    71 => x"7f3e0000",
    72 => x"7a7b4941",
    73 => x"7f7f0000",
    74 => x"7f7f0808",
    75 => x"41000000",
    76 => x"00417f7f",
    77 => x"60200000",
    78 => x"3f7f4040",
    79 => x"087f7f00",
    80 => x"4163361c",
    81 => x"7f7f0000",
    82 => x"40404040",
    83 => x"067f7f00",
    84 => x"7f7f060c",
    85 => x"067f7f00",
    86 => x"7f7f180c",
    87 => x"7f3e0000",
    88 => x"3e7f4141",
    89 => x"7f7f0000",
    90 => x"060f0909",
    91 => x"417f3e00",
    92 => x"407e7f61",
    93 => x"7f7f0000",
    94 => x"667f1909",
    95 => x"6f260000",
    96 => x"327b594d",
    97 => x"01010000",
    98 => x"01017f7f",
    99 => x"7f3f0000",
   100 => x"3f7f4040",
   101 => x"3f0f0000",
   102 => x"0f3f7070",
   103 => x"307f7f00",
   104 => x"7f7f3018",
   105 => x"36634100",
   106 => x"63361c1c",
   107 => x"06030141",
   108 => x"03067c7c",
   109 => x"59716101",
   110 => x"4143474d",
   111 => x"7f000000",
   112 => x"0041417f",
   113 => x"06030100",
   114 => x"6030180c",
   115 => x"41000040",
   116 => x"007f7f41",
   117 => x"060c0800",
   118 => x"080c0603",
   119 => x"80808000",
   120 => x"80808080",
   121 => x"00000000",
   122 => x"00040703",
   123 => x"74200000",
   124 => x"787c5454",
   125 => x"7f7f0000",
   126 => x"387c4444",
   127 => x"7c380000",
   128 => x"00444444",
   129 => x"7c380000",
   130 => x"7f7f4444",
   131 => x"7c380000",
   132 => x"185c5454",
   133 => x"7e040000",
   134 => x"0005057f",
   135 => x"bc180000",
   136 => x"7cfca4a4",
   137 => x"7f7f0000",
   138 => x"787c0404",
   139 => x"00000000",
   140 => x"00407d3d",
   141 => x"80800000",
   142 => x"007dfd80",
   143 => x"7f7f0000",
   144 => x"446c3810",
   145 => x"00000000",
   146 => x"00407f3f",
   147 => x"0c7c7c00",
   148 => x"787c0c18",
   149 => x"7c7c0000",
   150 => x"787c0404",
   151 => x"7c380000",
   152 => x"387c4444",
   153 => x"fcfc0000",
   154 => x"183c2424",
   155 => x"3c180000",
   156 => x"fcfc2424",
   157 => x"7c7c0000",
   158 => x"080c0404",
   159 => x"5c480000",
   160 => x"20745454",
   161 => x"3f040000",
   162 => x"0044447f",
   163 => x"7c3c0000",
   164 => x"7c7c4040",
   165 => x"3c1c0000",
   166 => x"1c3c6060",
   167 => x"607c3c00",
   168 => x"3c7c6030",
   169 => x"386c4400",
   170 => x"446c3810",
   171 => x"bc1c0000",
   172 => x"1c3c60e0",
   173 => x"64440000",
   174 => x"444c5c74",
   175 => x"08080000",
   176 => x"4141773e",
   177 => x"00000000",
   178 => x"00007f7f",
   179 => x"41410000",
   180 => x"08083e77",
   181 => x"01010200",
   182 => x"01020203",
   183 => x"7f7f7f00",
   184 => x"7f7f7f7f",
   185 => x"1c080800",
   186 => x"7f3e3e1c",
   187 => x"3e7f7f7f",
   188 => x"081c1c3e",
   189 => x"18100008",
   190 => x"10187c7c",
   191 => x"30100000",
   192 => x"10307c7c",
   193 => x"60301000",
   194 => x"061e7860",
   195 => x"3c664200",
   196 => x"42663c18",
   197 => x"6a387800",
   198 => x"386cc6c2",
   199 => x"00006000",
   200 => x"60000060",
   201 => x"5b5e0e00",
   202 => x"1e0e5d5c",
   203 => x"f9c24c71",
   204 => x"c04dbfe2",
   205 => x"741ec04b",
   206 => x"87c702ab",
   207 => x"c048a6c4",
   208 => x"c487c578",
   209 => x"78c148a6",
   210 => x"731e66c4",
   211 => x"87dfee49",
   212 => x"e0c086c8",
   213 => x"87efef49",
   214 => x"6a4aa5c4",
   215 => x"87f0f049",
   216 => x"cb87c6f1",
   217 => x"c883c185",
   218 => x"ff04abb7",
   219 => x"262687c7",
   220 => x"264c264d",
   221 => x"1e4f264b",
   222 => x"f9c24a71",
   223 => x"f9c25ae6",
   224 => x"78c748e6",
   225 => x"87ddfe49",
   226 => x"731e4f26",
   227 => x"c04a711e",
   228 => x"d303aab7",
   229 => x"eadbc287",
   230 => x"87c405bf",
   231 => x"87c24bc1",
   232 => x"dbc24bc0",
   233 => x"87c45bee",
   234 => x"5aeedbc2",
   235 => x"bfeadbc2",
   236 => x"c19ac14a",
   237 => x"ec49a2c0",
   238 => x"48fc87e8",
   239 => x"bfeadbc2",
   240 => x"87effe78",
   241 => x"c44a711e",
   242 => x"49721e66",
   243 => x"87dedfff",
   244 => x"1e4f2626",
   245 => x"bfeadbc2",
   246 => x"cedcff49",
   247 => x"daf9c287",
   248 => x"78bfe848",
   249 => x"48d6f9c2",
   250 => x"c278bfec",
   251 => x"4abfdaf9",
   252 => x"99ffc349",
   253 => x"722ab7c8",
   254 => x"c2b07148",
   255 => x"2658e2f9",
   256 => x"5b5e0e4f",
   257 => x"710e5d5c",
   258 => x"87c7ff4b",
   259 => x"48d5f9c2",
   260 => x"497350c0",
   261 => x"87f3dbff",
   262 => x"c24c4970",
   263 => x"49eecb9c",
   264 => x"7087cfcb",
   265 => x"f9c24d49",
   266 => x"05bf97d5",
   267 => x"d087e4c1",
   268 => x"f9c24966",
   269 => x"0599bfde",
   270 => x"66d487d7",
   271 => x"d6f9c249",
   272 => x"cc0599bf",
   273 => x"ff497387",
   274 => x"7087c0db",
   275 => x"c2c10298",
   276 => x"fd4cc187",
   277 => x"497587fd",
   278 => x"7087e3ca",
   279 => x"87c60298",
   280 => x"48d5f9c2",
   281 => x"f9c250c1",
   282 => x"05bf97d5",
   283 => x"c287e4c0",
   284 => x"49bfdef9",
   285 => x"059966d0",
   286 => x"c287d6ff",
   287 => x"49bfd6f9",
   288 => x"059966d4",
   289 => x"7387caff",
   290 => x"fed9ff49",
   291 => x"05987087",
   292 => x"7487fefe",
   293 => x"87d7fb48",
   294 => x"5c5b5e0e",
   295 => x"86f40e5d",
   296 => x"ec4c4dc0",
   297 => x"a6c47ebf",
   298 => x"e2f9c248",
   299 => x"1ec178bf",
   300 => x"49c71ec0",
   301 => x"c887cafd",
   302 => x"02987086",
   303 => x"49ff87ce",
   304 => x"c187c7fb",
   305 => x"d9ff49da",
   306 => x"4dc187c1",
   307 => x"97d5f9c2",
   308 => x"87c302bf",
   309 => x"c287f9cd",
   310 => x"4bbfdaf9",
   311 => x"bfeadbc2",
   312 => x"87ebc005",
   313 => x"ff49fdc3",
   314 => x"c387e0d8",
   315 => x"d8ff49fa",
   316 => x"497387d9",
   317 => x"7199ffc3",
   318 => x"fb49c01e",
   319 => x"497387c6",
   320 => x"7129b7c8",
   321 => x"fa49c11e",
   322 => x"86c887fa",
   323 => x"c287c1c6",
   324 => x"4bbfdef9",
   325 => x"87dd029b",
   326 => x"bfe6dbc2",
   327 => x"87dec749",
   328 => x"c4059870",
   329 => x"d24bc087",
   330 => x"49e0c287",
   331 => x"c287c3c7",
   332 => x"c658eadb",
   333 => x"e6dbc287",
   334 => x"7378c048",
   335 => x"0599c249",
   336 => x"ebc387ce",
   337 => x"c2d7ff49",
   338 => x"c2497087",
   339 => x"87c20299",
   340 => x"49734cfb",
   341 => x"ce0599c1",
   342 => x"49f4c387",
   343 => x"87ebd6ff",
   344 => x"99c24970",
   345 => x"fa87c202",
   346 => x"c849734c",
   347 => x"87ce0599",
   348 => x"ff49f5c3",
   349 => x"7087d4d6",
   350 => x"0299c249",
   351 => x"f9c287d5",
   352 => x"ca02bfe6",
   353 => x"88c14887",
   354 => x"58eaf9c2",
   355 => x"ff87c2c0",
   356 => x"734dc14c",
   357 => x"0599c449",
   358 => x"f2c387ce",
   359 => x"ead5ff49",
   360 => x"c2497087",
   361 => x"87dc0299",
   362 => x"bfe6f9c2",
   363 => x"b7c7487e",
   364 => x"cbc003a8",
   365 => x"c1486e87",
   366 => x"eaf9c280",
   367 => x"87c2c058",
   368 => x"4dc14cfe",
   369 => x"ff49fdc3",
   370 => x"7087c0d5",
   371 => x"0299c249",
   372 => x"c287d5c0",
   373 => x"02bfe6f9",
   374 => x"c287c9c0",
   375 => x"c048e6f9",
   376 => x"87c2c078",
   377 => x"4dc14cfd",
   378 => x"ff49fac3",
   379 => x"7087dcd4",
   380 => x"0299c249",
   381 => x"c287d9c0",
   382 => x"48bfe6f9",
   383 => x"03a8b7c7",
   384 => x"c287c9c0",
   385 => x"c748e6f9",
   386 => x"87c2c078",
   387 => x"4dc14cfc",
   388 => x"03acb7c0",
   389 => x"c487d1c0",
   390 => x"d8c14a66",
   391 => x"c0026a82",
   392 => x"4b6a87c6",
   393 => x"0f734974",
   394 => x"f0c31ec0",
   395 => x"49dac11e",
   396 => x"c887cef7",
   397 => x"02987086",
   398 => x"c887e2c0",
   399 => x"f9c248a6",
   400 => x"c878bfe6",
   401 => x"91cb4966",
   402 => x"714866c4",
   403 => x"6e7e7080",
   404 => x"c8c002bf",
   405 => x"4bbf6e87",
   406 => x"734966c8",
   407 => x"029d750f",
   408 => x"c287c8c0",
   409 => x"49bfe6f9",
   410 => x"c287faf2",
   411 => x"02bfeedb",
   412 => x"4987ddc0",
   413 => x"7087c7c2",
   414 => x"d3c00298",
   415 => x"e6f9c287",
   416 => x"e0f249bf",
   417 => x"f449c087",
   418 => x"dbc287c0",
   419 => x"78c048ee",
   420 => x"daf38ef4",
   421 => x"5b5e0e87",
   422 => x"1e0e5d5c",
   423 => x"f9c24c71",
   424 => x"c149bfe2",
   425 => x"c14da1cd",
   426 => x"7e6981d1",
   427 => x"cf029c74",
   428 => x"4ba5c487",
   429 => x"f9c27b74",
   430 => x"f249bfe2",
   431 => x"7b6e87f9",
   432 => x"c4059c74",
   433 => x"c24bc087",
   434 => x"734bc187",
   435 => x"87faf249",
   436 => x"c70266d4",
   437 => x"87da4987",
   438 => x"87c24a70",
   439 => x"dbc24ac0",
   440 => x"f2265af2",
   441 => x"000087c9",
   442 => x"00000000",
   443 => x"00000000",
   444 => x"711e0000",
   445 => x"bfc8ff4a",
   446 => x"48a17249",
   447 => x"ff1e4f26",
   448 => x"fe89bfc8",
   449 => x"c0c0c0c0",
   450 => x"c401a9c0",
   451 => x"c24ac087",
   452 => x"724ac187",
   453 => x"0e4f2648",
   454 => x"5d5c5b5e",
   455 => x"4d711e0e",
   456 => x"754bd4ff",
   457 => x"eaf9c21e",
   458 => x"c4c3fe49",
   459 => x"7086c487",
   460 => x"c3026e7e",
   461 => x"f9c287ff",
   462 => x"754cbff2",
   463 => x"f4ddfe49",
   464 => x"05a8de87",
   465 => x"7587ebc0",
   466 => x"ecd3ff49",
   467 => x"02987087",
   468 => x"f8c287db",
   469 => x"c01ebfed",
   470 => x"d0ff49e1",
   471 => x"86c487fb",
   472 => x"48cfe1c2",
   473 => x"f8c250c0",
   474 => x"eafe49f9",
   475 => x"c348c187",
   476 => x"d0ff87c5",
   477 => x"78c5c848",
   478 => x"c07bd6c1",
   479 => x"bf976e4a",
   480 => x"c1486e7b",
   481 => x"c17e7080",
   482 => x"b7e0c082",
   483 => x"ecff04aa",
   484 => x"48d0ff87",
   485 => x"c5c878c4",
   486 => x"7bd3c178",
   487 => x"78c47bc1",
   488 => x"c1029c74",
   489 => x"e7c287fd",
   490 => x"c0c87ee6",
   491 => x"b7c08c4d",
   492 => x"87c603ac",
   493 => x"4da4c0c8",
   494 => x"f4c24cc0",
   495 => x"49bf97d7",
   496 => x"d20299d0",
   497 => x"c21ec087",
   498 => x"fe49eaf9",
   499 => x"c487f7c3",
   500 => x"4a497086",
   501 => x"c287efc0",
   502 => x"c21ee6e7",
   503 => x"fe49eaf9",
   504 => x"c487e3c3",
   505 => x"4a497086",
   506 => x"c848d0ff",
   507 => x"d4c178c5",
   508 => x"bf976e7b",
   509 => x"c1486e7b",
   510 => x"c17e7080",
   511 => x"f0ff058d",
   512 => x"48d0ff87",
   513 => x"9a7278c4",
   514 => x"87c5c005",
   515 => x"e6c048c0",
   516 => x"c21ec187",
   517 => x"fe49eaf9",
   518 => x"c487d1c1",
   519 => x"059c7486",
   520 => x"ff87c3fe",
   521 => x"c5c848d0",
   522 => x"7bd3c178",
   523 => x"78c47bc0",
   524 => x"c2c048c1",
   525 => x"2648c087",
   526 => x"4c264d26",
   527 => x"4f264b26",
   528 => x"c44a711e",
   529 => x"87c50566",
   530 => x"cafb4972",
   531 => x"004f2687",
   532 => x"dee2c21e",
   533 => x"b9c149bf",
   534 => x"59e2e2c2",
   535 => x"c348d4ff",
   536 => x"d0ff78ff",
   537 => x"78e1c848",
   538 => x"c148d4ff",
   539 => x"7131c478",
   540 => x"48d0ff78",
   541 => x"2678e0c0",
   542 => x"e2c21e4f",
   543 => x"f9c21ed2",
   544 => x"fdfd49ea",
   545 => x"86c487eb",
   546 => x"c3029870",
   547 => x"87c0ff87",
   548 => x"35314f26",
   549 => x"205a484b",
   550 => x"46432020",
   551 => x"00000047",
   552 => x"5e0e0000",
   553 => x"0e5d5c5b",
   554 => x"bfd6f9c2",
   555 => x"cbe4c24a",
   556 => x"724c49bf",
   557 => x"ff4d71bc",
   558 => x"c087e6c1",
   559 => x"d049744b",
   560 => x"e7c00299",
   561 => x"48d0ff87",
   562 => x"ff78e1c8",
   563 => x"78c548d4",
   564 => x"99d04975",
   565 => x"c387c302",
   566 => x"e6c278f0",
   567 => x"817349f7",
   568 => x"d4ff4811",
   569 => x"d0ff7808",
   570 => x"78e0c048",
   571 => x"832d2cc1",
   572 => x"ff04abc8",
   573 => x"c0ff87c7",
   574 => x"e4c287df",
   575 => x"f9c248cb",
   576 => x"2678bfd6",
   577 => x"264c264d",
   578 => x"004f264b",
   579 => x"1e000000",
   580 => x"4bc01e73",
   581 => x"48cfe1c2",
   582 => x"1ec850de",
   583 => x"49fef9c2",
   584 => x"87d0d5fe",
   585 => x"1e7286c4",
   586 => x"48c0e6c2",
   587 => x"49c6fac2",
   588 => x"204aa1c4",
   589 => x"05aa7141",
   590 => x"4a2687f9",
   591 => x"49c4e6c2",
   592 => x"87cef9fd",
   593 => x"029a4a70",
   594 => x"fe4987c5",
   595 => x"7287efc7",
   596 => x"d0e6c21e",
   597 => x"c6fac248",
   598 => x"4aa1c449",
   599 => x"aa714120",
   600 => x"2687f905",
   601 => x"fef9c24a",
   602 => x"87ebf649",
   603 => x"c4059870",
   604 => x"d4e6c287",
   605 => x"fe49c04b",
   606 => x"7387e5c5",
   607 => x"87c7fe48",
   608 => x"00202020",
   609 => x"45544f4a",
   610 => x"20204f47",
   611 => x"00202020",
   612 => x"00435241",
   613 => x"20435241",
   614 => x"20746f6e",
   615 => x"6e756f66",
   616 => x"4c202e64",
   617 => x"2064616f",
   618 => x"00435241",
   619 => x"87e8eb1e",
   620 => x"f887effb",
   621 => x"164f2687",
   622 => x"2e25261e",
   623 => x"2e3e3d36",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
