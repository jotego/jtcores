localparam [1:0] SYS_INFO    = 2'b01,
                 TARGET_INFO = 2'b10;
