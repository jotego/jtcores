localparam [1:0] VULGUS=2'b1,
                 HIGEMARU=2'd2;
