localparam [12:1] FILL={SCR1,8'd0};

localparam [3:0] OBJ=0, TEXT=1, SCR1=2, SCR2=3;
localparam [4:0] SEL_TXT=1,SEL_SCR1=2,SEL_SCR2=4,SEL_OBJ=8,SEL_NONE=16;
localparam [2:0] REGISTER_FINAL_COLOR=6;