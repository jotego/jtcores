/*  This file is part of JTFRAME.
    JTFRAME program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTFRAME program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTFRAME.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 8-5-2021 */

// ctrl+shift selects sys info
// alt+shift selects target info

module jtframe_debug #(
    parameter COLORW=4
) (
    input              clk,
    input              rst,

    input              shift,         // count step 16, instead of 1
    input              ctrl,          // reset debug_bus
    input              alt,
    input              debug_plus,
    input              debug_minus,
    input              debug_rst,
    input        [3:0] key_gfx, board_gfx,
    input        [5:0] key_snd,               // enable individual sound channels
    input        [7:0] key_digit,
    // overlay the value on video
    input              pxl_cen,
    input [COLORW-1:0] rin,
    input [COLORW-1:0] gin,
    input [COLORW-1:0] bin,
    input              lhbl,
    input              lvbl,
    input              dip_flip,

    // combinational output
    output [COLORW-1:0] rout,
    output [COLORW-1:0] gout,
    output [COLORW-1:0] bout,
    // debug features
    output        [7:0] debug_bus,
    input         [7:0] debug_view, // an 8-bit signal that will be shown over the game image
    input         [7:0] sys_info,   // system information generated within JTFRAME, not the game
    input         [7:0] target_info,  // system information generated by the JTFRAME target, not the game
    input         [7:0] snd_vol,
    input               snd_mode,
    output        [3:0] gfx_en,
    output        [5:0] snd_en
);

reg  [2:0] color;
reg  [7:0] view_mux;
reg        vtoggle_l;
reg  [1:0] view_sel;
wire       vtoggle;

assign vtoggle = shift & ctrl;

localparam [1:0] SYS_INFO    = 2'b01,
                 TARGET_INFO = 2'b10;

always @(posedge clk) begin
    if( rst ) begin
        view_sel   <= 0;
        view_mux   <= 0;
    end else begin
        vtoggle_l  <= vtoggle;

        if( vtoggle && !vtoggle_l ) begin
            view_sel <= view_sel==2 ? 2'd0 : view_sel+1'd1;
        end
        case( view_sel )
            default:     view_mux <= debug_view;
            SYS_INFO:    view_mux <= sys_info;
            TARGET_INFO: view_mux <= target_info;
        endcase
    end
end

// Video overlay
localparam [8:0] JTFRAME_DEBUG_VPOS=`JTFRAME_DEBUG_VPOS;

reg  [7:0] dmux;
wire [8:0] HBIN=((`JTFRAME_WIDTH&9'h1f8)>>1)-9'h10,
                 HHEX=HBIN+9'h44,
                 VOSD=(`JTFRAME_HEIGHT & 9'h1f8)-9'd8*JTFRAME_DEBUG_VPOS, // 4 rows above bottom
                 VVIEW=VOSD+9'd8*9'd2;

wire [8:0] veff, heff;
wire       osd_on = debug_view_sel | debug_bus_sel;
reg        debug_view_sel, debug_bus_sel, hex_col, bin_col, hex_en, bin_en;

always @(posedge clk) begin
    color <= 7;
    if( view_sel==SYS_INFO    ) color<=3'b100; // system info is shown reddish
    if( view_sel==TARGET_INFO ) color<=3'b001; // system info is shown blueish
end

always @(posedge clk) begin
    // display of debug_bus
    debug_bus_sel  <=  debug_bus!=0 && veff[8:3]==VOSD[8:3];
    debug_view_sel <= (view_mux !=0 || view_sel!=0 || debug_bus!=0) && veff[8:3]==VVIEW[8:3];

    hex_col <= heff[8:4] == HHEX[8:4];
    bin_col <= heff[8:6] == HBIN[8:6];
    if(pxl_cen) begin
        hex_en <= osd_on & hex_col;
        bin_en <= osd_on & bin_col;
        dmux   <= debug_view_sel ? view_mux : debug_bus;
    end
end

wire [3:0] gfx_toggle = key_gfx | board_gfx;

jtframe_toggle #(.W(4),.VALUE_AT_RST(1'b1)) u_gfxen(
    .rst        ( rst         ),
    .clk        ( clk         ),
    .toggle     ( gfx_toggle  ),
    .q          ( gfx_en      )
);

jtframe_toggle #(.W(6),.VALUE_AT_RST(1'b1)) u_snd(
    .rst        ( rst         ),
    .clk        ( clk         ),
    .toggle     ( key_snd     ),
    .q          ( snd_en      )
);

jtframe_binhex_overlay #(.COLORW(COLORW)) u_overlay(
    .clk        ( clk         ),
    .v          ( veff        ),
    .h          ( heff        ),

    .bin_en     ( bin_en      ),
    .hex_en     ( hex_en      ),
    .din        ( dmux        ),
    .color      ( color       ),

    .rin        ( rin         ),
    .gin        ( gin         ),
    .bin        ( bin         ),

    .rout       ( rout        ),
    .gout       ( gout        ),
    .bout       ( bout        )
);

jtframe_video_counter u_vcounters(
    .rst        ( rst         ),
    .clk        ( clk         ),
    .pxl_cen    ( pxl_cen     ),

    .lhbl       ( lhbl        ),
    .lvbl       ( lvbl        ),
    .flip       ( dip_flip    ),

    .v          ( veff        ),
    .h          ( heff        )
);

jtframe_debug_bus u_debug_bus(
    .rst        ( rst         ),
    .clk        ( clk         ),
    .shift      ( shift       ),
    .ctrl       ( ctrl        ),
    .inc        ( debug_plus  ),
    .dec        ( debug_minus ),
    .key_digit  ( key_digit   ),
    .debug_bus  ( debug_bus   )
);

endmodule