../../shouse/hdl/vtimer.vh