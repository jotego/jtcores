/*  This file is part of JTCORES.
    JTCORES program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTCORES program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTCORES.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 3-4-2022 */

module jtrastan_snd(
    input                rst,
    input                clk,
    input                cen4, cen2, cen_pcm,

    // From main CPU
    input                main_addr,
    input         [ 3:0] main_dout,
    output        [ 3:0] main_din,
    input                main_rnw,
    input                sn_rd,
    input                sn_we,

    output        [15:0] rom_addr,
    output reg           rom_cs,
    input                rom_ok,
    input         [ 7:0] rom_data,

    output reg    [15:0] pcm_addr,
    output reg           pcm_cs,
    input                pcm_ok,
    input         [ 7:0] pcm_data,

    output signed [15:0] fm_l, fm_r,
    output signed [11:0] pcm
);
`ifndef NOSOUND
wire signed [15:0] pre_snd, left_opm, right_opm;
wire signed [11:0] pcm_snd;
wire               int_n, rfsh_n;
wire        [15:0] A;
wire        [ 7:0] dout, opm_dout, ram_dout;
wire        [ 3:0] pc6_dout;
reg                opm_cs, opl_cs, ram_cs, pc6_cs;
reg                pcm_rst, pcm_stop, pcm_start, pcm_addr_cs;
wire               rd_n, wr_n, mreq_n, nmi_n;
wire               ct1, ct2, vclk, pc6_rst, mem_acc;
reg                nibble_sel, vclk_l, snd_rstn;
reg         [15:0] pcm_cnt;
wire        [ 3:0] pcm_nibble;
reg         [ 7:0] din;
wire               pc60_rd, pc60_we;

assign mem_acc    = rfsh_n && !mreq_n;
assign rom_addr   = A[14] ? { ct2, ct1, A[13:0]  } : A;
assign pcm_nibble = !nibble_sel ? pcm_data[7:4] : pcm_data[3:0];
assign pc60_rd    = pc6_cs && !rd_n;
assign pc60_we    = pc6_cs && !wr_n;

always @(posedge clk) begin
    snd_rstn <= ~(rst | pc6_rst);
end

// PCM controller
always @(posedge clk) begin
    if( rst ) begin
        pcm_addr   <= 0;
        pcm_cs     <= 0;
        nibble_sel <= 0;
        pcm_rst    <= 1;
    end else begin
        vclk_l <= vclk;
        if( pcm_addr_cs ) pcm_addr[15:8] <= dout;
        if( pcm_start ) begin
            pcm_cs         <= 1;
            pcm_rst        <= 0;
            pcm_addr[ 7:0] <= 0;
            nibble_sel     <= 0;
        end
        if( pcm_stop    ) begin
            pcm_cs         <= 0;
            pcm_rst        <= 1;
        end
        if( vclk && ! vclk_l && !pcm_rst)
            { pcm_addr, nibble_sel } <= { pcm_addr, nibble_sel } + 1'd1;
    end
end

always @* begin
    rom_cs      = !A[15] && !rd_n && mem_acc;
    ram_cs      = 0;
    opm_cs      = 0;
    pc6_cs      = 0;
    pcm_addr_cs = 0;
    pcm_start   = 0;
    pcm_stop    = 0;
    if( mem_acc && A[15]) begin
        case( A[14:12] )
            0: ram_cs = 1;
            1: opm_cs = 1;
            2: pc6_cs = 1;
            3: pcm_addr_cs = !wr_n;
            4: pcm_start   = !wr_n;
            5: pcm_stop    = !wr_n;
            default:;
        endcase
    end
end

always @(posedge clk) begin
    din <=  rom_cs ? rom_data :
            ram_cs ? ram_dout :
            opm_cs ? opm_dout :
            pc6_cs ? { 4'hf, pc6_dout } :
                     8'h00;
end

jtrastan_pc060 u_pc060(
    .rst        ( rst       ),
    .clk        ( clk       ),

    .main_dout  ( main_dout ),
    .main_din   ( main_din  ),
    .main_addr  ( main_addr ),
    .main_rd    ( sn_rd     ),
    .main_we    ( sn_we     ),

    .snd_dout   ( dout[3:0] ),
    .snd_din    ( pc6_dout  ),
    .snd_addr   ( A[0]      ),
    .snd_rd     ( pc60_rd   ),
    .snd_we     ( pc60_we   ),
    .snd_nmin   ( nmi_n     ),
    .snd_rst    ( pc6_rst   )
);

jtframe_sysz80 u_cpu(
    .rst_n      ( snd_rstn  ),
    .clk        ( clk       ),
    .cen        ( cen4      ),
    .cpu_cen    (           ),
    .int_n      ( int_n     ),
    .nmi_n      ( nmi_n     ),
    .busrq_n    ( 1'b1      ),
    .m1_n       (           ),
    .mreq_n     ( mreq_n    ),
    .iorq_n     (           ),
    .rd_n       ( rd_n      ),
    .wr_n       ( wr_n      ),
    .rfsh_n     ( rfsh_n    ),
    .halt_n     (           ),
    .busak_n    (           ),
    .A          ( A         ),
    .cpu_din    ( din       ),
    .cpu_dout   ( dout      ),
    .ram_dout   ( ram_dout  ),
    // ROM access
    .ram_cs     ( ram_cs    ),
    .rom_cs     ( rom_cs    ),
    .rom_ok     ( rom_ok    )
);

jt51 u_jt51(
    .rst    ( ~snd_rstn ),
    .clk    ( clk       ),
    .cen    ( cen4      ),
    .cen_p1 ( cen2      ),
    .cs_n   ( ~opm_cs   ),
    .wr_n   ( wr_n      ),
    .a0     ( A[0]       ),
    .din    ( dout      ),
    .dout   ( opm_dout  ),
    // peripheral control
    .ct1    ( ct1       ),
    .ct2    ( ct2       ),
    .irq_n  ( int_n     ),
    // Low resolution output (same as real chip)
    .sample (           ),
    .left   (           ),
    .right  (           ),
    // Full resolution output
    .xleft  ( fm_l      ),
    .xright ( fm_r      )
);

jt5205 u_5205( // 8kHz, 4 bits/sample
    .rst    ( pcm_rst   ),
    .clk    ( clk       ),
    .cen    ( cen_pcm   ),
    .sel    ( 2'b10     ),
    .din    ( pcm_nibble),
    .sound  ( pcm       ),
    .sample (           ),
    .irq    (           ),
    .vclk_o ( vclk      )
);
`else
assign main_din=0, rom_addr=0, fm_l=0, fm_r=0, pcm=0;
initial begin
    rom_cs=0;
    pcm_addr=0;
    pcm_cs=0;
end
`endif
endmodule
